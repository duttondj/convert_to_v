/////////////////////////////////////////////////////////////////////////////
//
// FILENAME: character_rom.v
//
// CREATED BY: <various online sources, fancy editing>
//
// DESCRIPTION: 
//    The appearance of the characters on the screen is determined by a "font 
//    ROM". The font ROM contains the pattern of pixels that should be 
//    displayed on the screen when a particular character needs to be 
//    displayed. The bits within the font ROM indicate which pixels of a 
//    8 x 16 bit tile should be displayed in the 'foreground' and which 
//    pixels on the display should be displayed in the background. A '1' 
//    in the font ROM indicates the corresponding pixel should be displayed 
//    in the foreground (i.e., white in our case) while a '0' in the font 
//    ROM indicates that the corresponding pixel should be blanked or put 
//    in the background (black in our case).
//
/////////////////////////////////////////////////////////////////////////////

module character_rom ( input clk, input [10:0] addr, output reg [7:0] rom);
	always@(posedge clk) begin
	   case(addr)
    // code x00
            11'd0:      rom = 8'b00000000;    // 0
            11'd1:      rom = 8'b00000000;    // 1
            11'd2:      rom = 8'b00000000;    // 2
            11'd3:      rom = 8'b00000000;    // 3
            11'd4:      rom = 8'b00000000;    // 4
            11'd5:      rom = 8'b00000000;    // 5
            11'd6:      rom = 8'b00000000;    // 6
            11'd7:      rom = 8'b00000000;    // 7
            11'd8:      rom = 8'b00000000;    // 8
            11'd9:      rom = 8'b00000000;    // 9
            11'd10:     rom = 8'b00000000;    // a
            11'd11:     rom = 8'b00000000;    // b
            11'd12:     rom = 8'b00000000;    // c
            11'd13:     rom = 8'b00000000;    // d
            11'd14:     rom = 8'b00000000;    // e
            11'd15:     rom = 8'b00000000;    // f
   // code x0 1       
            11'd16:     rom = 8'b00000000;    // 0
            11'd17:     rom = 8'b00000000;    // 1
            11'd18:     rom = 8'b01111110;    // 2  ******
            11'd19:     rom = 8'b10000001;    // 3 *      *
            11'd20:     rom = 8'b10100101;    // 4 * *  * *
            11'd21:     rom = 8'b10000001;    // 5 *      *
            11'd22:     rom = 8'b10000001;    // 6 *      *
            11'd23:     rom = 8'b10111101;    // 7 * **** *
            11'd24:     rom = 8'b10011001;    // 8 *  **  *
            11'd25:     rom = 8'b10000001;    // 9 *      *
            11'd26:     rom = 8'b10000001;    // a *      *
            11'd27:     rom = 8'b01111110;    // b  ******
            11'd28:     rom = 8'b00000000;    // c
            11'd29:     rom = 8'b00000000;    // d
            11'd30:     rom = 8'b00000000;    // e
            11'd31:     rom = 8'b00000000;    // f
   // code x02        
            11'd32:     rom = 8'b00000000;    // 0
            11'd33:     rom = 8'b00000000;    // 1
            11'd34:     rom = 8'b01111110;    // 2  ******
            11'd35:     rom = 8'b11111111;    // 3 ********
            11'd36:     rom = 8'b11011011;    // 4 ** ** **
            11'd37:     rom = 8'b11111111;    // 5 ********
            11'd38:     rom = 8'b11111111;    // 6 ********
            11'd39:     rom = 8'b11000011;    // 7 **    **
            11'd40:     rom = 8'b11100111;    // 8 ***  ***
            11'd41:     rom = 8'b11111111;    // 9 ********
            11'd42:     rom = 8'b11111111;    // a ********
            11'd43:     rom = 8'b01111110;    // b  ******
            11'd44:     rom = 8'b00000000;    // c
            11'd45:     rom = 8'b00000000;    // d
            11'd46:     rom = 8'b00000000;    // e
            11'd47:     rom = 8'b00000000;    // f
   // code x03        
            11'd48:     rom = 8'b00000000;    // 0
            11'd49:     rom = 8'b00000000;    // 1
            11'd50:     rom = 8'b00000000;    // 2
            11'd51:     rom = 8'b00000000;    // 3
            11'd52:     rom = 8'b01101100;    // 4  ** **
            11'd53:     rom = 8'b11111110;    // 5 *******
            11'd54:     rom = 8'b11111110;    // 6 *******
            11'd55:     rom = 8'b11111110;    // 7 *******
            11'd56:     rom = 8'b11111110;    // 8 *******
            11'd57:     rom = 8'b01111100;    // 9  *****
            11'd58:     rom = 8'b00111000;    // a   ***
            11'd59:     rom = 8'b00010000;    // b    *
            11'd60:     rom = 8'b00000000;    // c
            11'd61:     rom = 8'b00000000;    // d
            11'd62:     rom = 8'b00000000;    // e
            11'd63:     rom = 8'b00000000;    // f
   // code x04        
            11'd64:     rom = 8'b00000000;    // 0
            11'd65:     rom = 8'b00000000;    // 1
            11'd66:     rom = 8'b00000000;    // 2
            11'd67:     rom = 8'b00000000;    // 3
            11'd68:     rom = 8'b00010000;    // 4    *
            11'd69:     rom = 8'b00111000;    // 5   ***
            11'd70:     rom = 8'b01111100;    // 6  *****
            11'd71:     rom = 8'b11111110;    // 7 *******
            11'd72:     rom = 8'b01111100;    // 8  *****
            11'd73:     rom = 8'b00111000;    // 9   ***
            11'd74:     rom = 8'b00010000;    // a    *
            11'd75:     rom = 8'b00000000;    // b
            11'd76:     rom = 8'b00000000;    // c
            11'd77:     rom = 8'b00000000;    // d
            11'd78:     rom = 8'b00000000;    // e
            11'd79:     rom = 8'b00000000;    // f
   // code x05        
            11'd80:     rom = 8'b00000000;    // 0
            11'd81:     rom = 8'b00000000;    // 1
            11'd82:     rom = 8'b00000000;    // 2
            11'd83:     rom = 8'b00011000;    // 3    **
            11'd84:     rom = 8'b00111100;    // 4   ****
            11'd85:     rom = 8'b00111100;    // 5   ****
            11'd86:     rom = 8'b11100111;    // 6 ***  ***
            11'd87:     rom = 8'b11100111;    // 7 ***  ***
            11'd88:     rom = 8'b11100111;    // 8 ***  ***
            11'd89:     rom = 8'b00011000;    // 9    **
            11'd90:     rom = 8'b00011000;    // a    **
            11'd91:     rom = 8'b00111100;    // b   ****
            11'd92:     rom = 8'b00000000;    // c
            11'd93:     rom = 8'b00000000;    // d
            11'd94:     rom = 8'b00000000;    // e
            11'd95:     rom = 8'b00000000;    // f
   // code x06        
            11'd96:     rom = 8'b00000000;    // 0
            11'd97:     rom = 8'b00000000;    // 1
            11'd98:     rom = 8'b00000000;    // 2
            11'd99:     rom = 8'b00011000;    // 3    **
            11'd100:    rom = 8'b00111100;    // 4   ****
            11'd101:    rom = 8'b01111110;    // 5  ******
            11'd102:    rom = 8'b11111111;    // 6 ********
            11'd103:    rom = 8'b11111111;    // 7 ********
            11'd104:    rom = 8'b01111110;    // 8  ******
            11'd105:    rom = 8'b00011000;    // 9    **
            11'd106:    rom = 8'b00011000;    // a    **
            11'd107:    rom = 8'b00111100;    // b   ****
            11'd108:    rom = 8'b00000000;    // c
            11'd109:    rom = 8'b00000000;    // d
            11'd110:    rom = 8'b00000000;    // e
            11'd111:    rom = 8'b00000000;    // f
   // code x07         
            11'd112:    rom = 8'b00000000;    // 0
            11'd113:    rom = 8'b00000000;    // 1
            11'd114:    rom = 8'b00000000;    // 2
            11'd115:    rom = 8'b00000000;    // 3
            11'd116:    rom = 8'b00000000;    // 4
            11'd117:    rom = 8'b00000000;    // 5
            11'd118:    rom = 8'b00011000;    // 6    **
            11'd119:    rom = 8'b00111100;    // 7   ****
            11'd120:    rom = 8'b00111100;    // 8   ****
            11'd121:    rom = 8'b00011000;    // 9    **
            11'd122:    rom = 8'b00000000;    // a
            11'd123:    rom = 8'b00000000;    // b
            11'd124:    rom = 8'b00000000;    // c
            11'd125:    rom = 8'b00000000;    // d
            11'd126:    rom = 8'b00000000;    // e
            11'd127:    rom = 8'b00000000;    // f
   // code x08         
            11'd128:    rom = 8'b11111111;    // 0 ********
            11'd129:    rom = 8'b11111111;    // 1 ********
            11'd130:    rom = 8'b11111111;    // 2 ********
            11'd131:    rom = 8'b11111111;    // 3 ********
            11'd132:    rom = 8'b11111111;    // 4 ********
            11'd133:    rom = 8'b11111111;    // 5 ********
            11'd134:    rom = 8'b11100111;    // 6 ***  ***
            11'd135:    rom = 8'b11000011;    // 7 **    **
            11'd136:    rom = 8'b11000011;    // 8 **    **
            11'd137:    rom = 8'b11100111;    // 9 ***  ***
            11'd138:    rom = 8'b11111111;    // a ********
            11'd139:    rom = 8'b11111111;    // b ********
            11'd140:    rom = 8'b11111111;    // c ********
            11'd141:    rom = 8'b11111111;    // d ********
            11'd142:    rom = 8'b11111111;    // e ********
            11'd143:    rom = 8'b11111111;    // f ********
   // code x09         
            11'd144:    rom = 8'b00000000;    // 0
            11'd145:    rom = 8'b00000000;    // 1
            11'd146:    rom = 8'b00000000;    // 2
            11'd147:    rom = 8'b00000000;    // 3
            11'd148:    rom = 8'b00000000;    // 4
            11'd149:    rom = 8'b00111100;    // 5   ****
            11'd150:    rom = 8'b01100110;    // 6  **  **
            11'd151:    rom = 8'b01000010;    // 7  *    *
            11'd152:    rom = 8'b01000010;    // 8  *    *
            11'd153:    rom = 8'b01100110;    // 9  **  **
            11'd154:    rom = 8'b00111100;    // a   ****
            11'd155:    rom = 8'b00000000;    // b
            11'd156:    rom = 8'b00000000;    // c
            11'd157:    rom = 8'b00000000;    // d
            11'd158:    rom = 8'b00000000;    // e
            11'd159:    rom = 8'b00000000;    // f
   // code x0a         
            11'd160:    rom = 8'b11111111;    // 0 ********
            11'd161:    rom = 8'b11111111;    // 1 ********
            11'd162:    rom = 8'b11111111;    // 2 ********
            11'd163:    rom = 8'b11111111;    // 3 ********
            11'd164:    rom = 8'b11111111;    // 4 ********
            11'd165:    rom = 8'b11000011;    // 5 **    **
            11'd166:    rom = 8'b10011001;    // 6 *  **  *
            11'd167:    rom = 8'b10111101;    // 7 * **** *
            11'd168:    rom = 8'b10111101;    // 8 * **** *
            11'd169:    rom = 8'b10011001;    // 9 *  **  *
            11'd170:    rom = 8'b11000011;    // a **    **
            11'd171:    rom = 8'b11111111;    // b ********
            11'd172:    rom = 8'b11111111;    // c ********
            11'd173:    rom = 8'b11111111;    // d ********
            11'd174:    rom = 8'b11111111;    // e ********
            11'd175:    rom = 8'b11111111;    // f ********
   // code x0b         
            11'd176:    rom = 8'b00000000;    // 0
            11'd177:    rom = 8'b00000000;    // 1
            11'd178:    rom = 8'b00011110;    // 2    ****
            11'd179:    rom = 8'b00001110;    // 3     ***
            11'd180:    rom = 8'b00011010;    // 4    ** *
            11'd181:    rom = 8'b00110010;    // 5   **  *
            11'd182:    rom = 8'b01111000;    // 6  ****
            11'd183:    rom = 8'b11001100;    // 7 **  **
            11'd184:    rom = 8'b11001100;    // 8 **  **
            11'd185:    rom = 8'b11001100;    // 9 **  **
            11'd186:    rom = 8'b11001100;    // a **  **
            11'd187:    rom = 8'b01111000;    // b  ****
            11'd188:    rom = 8'b00000000;    // c
            11'd189:    rom = 8'b00000000;    // d
            11'd190:    rom = 8'b00000000;    // e
            11'd191:    rom = 8'b00000000;    // f
   // code x0c         
            11'd192:    rom = 8'b00000000;    // 0
            11'd193:    rom = 8'b00000000;    // 1
            11'd194:    rom = 8'b00111100;    // 2   ****
            11'd195:    rom = 8'b01100110;    // 3  **  **
            11'd196:    rom = 8'b01100110;    // 4  **  **
            11'd197:    rom = 8'b01100110;    // 5  **  **
            11'd198:    rom = 8'b01100110;    // 6  **  **
            11'd199:    rom = 8'b00111100;    // 7   ****
            11'd200:    rom = 8'b00011000;    // 8    **
            11'd201:    rom = 8'b01111110;    // 9  ******
            11'd202:    rom = 8'b00011000;    // a    **
            11'd203:    rom = 8'b00011000;    // b    **
            11'd204:    rom = 8'b00000000;    // c
            11'd205:    rom = 8'b00000000;    // d
            11'd206:    rom = 8'b00000000;    // e
            11'd207:    rom = 8'b00000000;    // f
   // code x0d         
            11'd208:    rom = 8'b00000000;    // 0
            11'd209:    rom = 8'b00000000;    // 1
            11'd210:    rom = 8'b00111111;    // 2   ******
            11'd211:    rom = 8'b00110011;    // 3   **  **
            11'd212:    rom = 8'b00111111;    // 4   ******
            11'd213:    rom = 8'b00110000;    // 5   **
            11'd214:    rom = 8'b00110000;    // 6   **
            11'd215:    rom = 8'b00110000;    // 7   **
            11'd216:    rom = 8'b00110000;    // 8   **
            11'd217:    rom = 8'b01110000;    // 9  ***
            11'd218:    rom = 8'b11110000;    // a ****
            11'd219:    rom = 8'b11100000;    // b ***
            11'd220:    rom = 8'b00000000;    // c
            11'd221:    rom = 8'b00000000;    // d
            11'd222:    rom = 8'b00000000;    // e
            11'd223:    rom = 8'b00000000;    // f
   // code x0e         
            11'd224:    rom = 8'b00000000;    // 0
            11'd225:    rom = 8'b00000000;    // 1
            11'd226:    rom = 8'b01111111;    // 2  *******
            11'd227:    rom = 8'b01100011;    // 3  **   **
            11'd228:    rom = 8'b01111111;    // 4  *******
            11'd229:    rom = 8'b01100011;    // 5  **   **
            11'd230:    rom = 8'b01100011;    // 6  **   **
            11'd231:    rom = 8'b01100011;    // 7  **   **
            11'd232:    rom = 8'b01100011;    // 8  **   **
            11'd233:    rom = 8'b01100111;    // 9  **  ***
            11'd234:    rom = 8'b11100111;    // a ***  ***
            11'd235:    rom = 8'b11100110;    // b ***  **
            11'd236:    rom = 8'b11000000;    // c **
            11'd237:    rom = 8'b00000000;    // d
            11'd238:    rom = 8'b00000000;    // e
            11'd239:    rom = 8'b00000000;    // f
   // code x0f         
            11'd240:    rom = 8'b00000000;    // 0
            11'd241:    rom = 8'b00000000;    // 1
            11'd242:    rom = 8'b00000000;    // 2
            11'd243:    rom = 8'b00011000;    // 3    **
            11'd244:    rom = 8'b00011000;    // 4    **
            11'd245:    rom = 8'b11011011;    // 5 ** ** **
            11'd246:    rom = 8'b00111100;    // 6   ****
            11'd247:    rom = 8'b11100111;    // 7 ***  ***
            11'd248:    rom = 8'b00111100;    // 8   ****
            11'd249:    rom = 8'b11011011;    // 9 ** ** **
            11'd250:    rom = 8'b00011000;    // a    **
            11'd251:    rom = 8'b00011000;    // b    **
            11'd252:    rom = 8'b00000000;    // c
            11'd253:    rom = 8'b00000000;    // d
            11'd254:    rom = 8'b00000000;    // e
            11'd255:    rom = 8'b00000000;    // f
   // code x10         
            11'd256:    rom = 8'b00000000;    // 0
            11'd257:    rom = 8'b10000000;    // 1 *
            11'd258:    rom = 8'b11000000;    // 2 **
            11'd259:    rom = 8'b11100000;    // 3 ***
            11'd260:    rom = 8'b11110000;    // 4 ****
            11'd261:    rom = 8'b11111000;    // 5 *****
            11'd262:    rom = 8'b11111110;    // 6 *******
            11'd263:    rom = 8'b11111000;    // 7 *****
            11'd264:    rom = 8'b11110000;    // 8 ****
            11'd265:    rom = 8'b11100000;    // 9 ***
            11'd266:    rom = 8'b11000000;    // a **
            11'd267:    rom = 8'b10000000;    // b *
            11'd268:    rom = 8'b00000000;    // c
            11'd269:    rom = 8'b00000000;    // d
            11'd270:    rom = 8'b00000000;    // e
            11'd271:    rom = 8'b00000000;    // f
   // code x11         
            11'd272:    rom = 8'b00000000;    // 0
            11'd273:    rom = 8'b00000010;    // 1       *
            11'd274:    rom = 8'b00000110;    // 2      **
            11'd275:    rom = 8'b00001110;    // 3     ***
            11'd276:    rom = 8'b00011110;    // 4    ****
            11'd277:    rom = 8'b00111110;    // 5   *****
            11'd278:    rom = 8'b11111110;    // 6 *******
            11'd279:    rom = 8'b00111110;    // 7   *****
            11'd280:    rom = 8'b00011110;    // 8    ****
            11'd281:    rom = 8'b00001110;    // 9     ***
            11'd282:    rom = 8'b00000110;    // a      **
            11'd283:    rom = 8'b00000010;    // b       *
            11'd284:    rom = 8'b00000000;    // c
            11'd285:    rom = 8'b00000000;    // d
            11'd286:    rom = 8'b00000000;    // e
            11'd287:    rom = 8'b00000000;    // f
   // code x12         
            11'd288:    rom = 8'b00000000;    // 0
            11'd289:    rom = 8'b00000000;    // 1
            11'd290:    rom = 8'b00011000;    // 2    **
            11'd291:    rom = 8'b00111100;    // 3   ****
            11'd292:    rom = 8'b01111110;    // 4  ******
            11'd293:    rom = 8'b00011000;    // 5    **
            11'd294:    rom = 8'b00011000;    // 6    **
            11'd295:    rom = 8'b00011000;    // 7    **
            11'd296:    rom = 8'b01111110;    // 8  ******
            11'd297:    rom = 8'b00111100;    // 9   ****
            11'd298:    rom = 8'b00011000;    // a    **
            11'd299:    rom = 8'b00000000;    // b
            11'd300:    rom = 8'b00000000;    // c
            11'd301:    rom = 8'b00000000;    // d
            11'd302:    rom = 8'b00000000;    // e
            11'd303:    rom = 8'b00000000;    // f
   // code x13         
            11'd304:    rom = 8'b00000000;    // 0
            11'd305:    rom = 8'b00000000;    // 1
            11'd306:    rom = 8'b01100110;    // 2  **  **
            11'd307:    rom = 8'b01100110;    // 3  **  **
            11'd308:    rom = 8'b01100110;    // 4  **  **
            11'd309:    rom = 8'b01100110;    // 5  **  **
            11'd310:    rom = 8'b01100110;    // 6  **  **
            11'd311:    rom = 8'b01100110;    // 7  **  **
            11'd312:    rom = 8'b01100110;    // 8  **  **
            11'd313:    rom = 8'b00000000;    // 9
            11'd314:    rom = 8'b01100110;    // a  **  **
            11'd315:    rom = 8'b01100110;    // b  **  **
            11'd316:    rom = 8'b00000000;    // c
            11'd317:    rom = 8'b00000000;    // d
            11'd318:    rom = 8'b00000000;    // e
            11'd319:    rom = 8'b00000000;    // f
   // code x14         
            11'd320:    rom = 8'b00000000;    // 0
            11'd321:    rom = 8'b00000000;    // 1
            11'd322:    rom = 8'b01111111;    // 2  *******
            11'd323:    rom = 8'b11011011;    // 3 ** ** **
            11'd324:    rom = 8'b11011011;    // 4 ** ** **
            11'd325:    rom = 8'b11011011;    // 5 ** ** **
            11'd326:    rom = 8'b01111011;    // 6  **** **
            11'd327:    rom = 8'b00011011;    // 7    ** **
            11'd328:    rom = 8'b00011011;    // 8    ** **
            11'd329:    rom = 8'b00011011;    // 9    ** **
            11'd330:    rom = 8'b00011011;    // a    ** **
            11'd331:    rom = 8'b00011011;    // b    ** **
            11'd332:    rom = 8'b00000000;    // c
            11'd333:    rom = 8'b00000000;    // d
            11'd334:    rom = 8'b00000000;    // e
            11'd335:    rom = 8'b00000000;    // f
   // code x15         
            11'd336:    rom = 8'b00000000;    // 0
            11'd337:    rom = 8'b01111100;    // 1  *****
            11'd338:    rom = 8'b11000110;    // 2 **   **
            11'd339:    rom = 8'b01100000;    // 3  **
            11'd340:    rom = 8'b00111000;    // 4   ***
            11'd341:    rom = 8'b01101100;    // 5  ** **
            11'd342:    rom = 8'b11000110;    // 6 **   **
            11'd343:    rom = 8'b11000110;    // 7 **   **
            11'd344:    rom = 8'b01101100;    // 8  ** **
            11'd345:    rom = 8'b00111000;    // 9   ***
            11'd346:    rom = 8'b00001100;    // a     **
            11'd347:    rom = 8'b11000110;    // b **   **
            11'd348:    rom = 8'b01111100;    // c  *****
            11'd349:    rom = 8'b00000000;    // d
            11'd350:    rom = 8'b00000000;    // e
            11'd351:    rom = 8'b00000000;    // f
   // code x16         
            11'd352:    rom = 8'b00000000;    // 0
            11'd353:    rom = 8'b00000000;    // 1
            11'd354:    rom = 8'b00000000;    // 2
            11'd355:    rom = 8'b00000000;    // 3
            11'd356:    rom = 8'b00000000;    // 4
            11'd357:    rom = 8'b00000000;    // 5
            11'd358:    rom = 8'b00000000;    // 6
            11'd359:    rom = 8'b00000000;    // 7
            11'd360:    rom = 8'b11111110;    // 8 *******
            11'd361:    rom = 8'b11111110;    // 9 *******
            11'd362:    rom = 8'b11111110;    // a *******
            11'd363:    rom = 8'b11111110;    // b *******
            11'd364:    rom = 8'b00000000;    // c
            11'd365:    rom = 8'b00000000;    // d
            11'd366:    rom = 8'b00000000;    // e
            11'd367:    rom = 8'b00000000;    // f
   // code x17         
            11'd368:    rom = 8'b00000000;    // 0
            11'd369:    rom = 8'b00000000;    // 1
            11'd370:    rom = 8'b00011000;    // 2    **
            11'd371:    rom = 8'b00111100;    // 3   ****
            11'd372:    rom = 8'b01111110;    // 4  ******
            11'd373:    rom = 8'b00011000;    // 5    **
            11'd374:    rom = 8'b00011000;    // 6    **
            11'd375:    rom = 8'b00011000;    // 7    **
            11'd376:    rom = 8'b01111110;    // 8  ******
            11'd377:    rom = 8'b00111100;    // 9   ****
            11'd378:    rom = 8'b00011000;    // a    **
            11'd379:    rom = 8'b01111110;    // b  ******
            11'd380:    rom = 8'b00110000;    // c
            11'd381:    rom = 8'b00000000;    // d
            11'd382:    rom = 8'b00000000;    // e
            11'd383:    rom = 8'b00000000;    // f
   // code x18         
            11'd384:    rom = 8'b00000000;    // 0
            11'd385:    rom = 8'b00000000;    // 1
            11'd386:    rom = 8'b00011000;    // 2    **
            11'd387:    rom = 8'b00111100;    // 3   ****
            11'd388:    rom = 8'b01111110;    // 4  ******
            11'd389:    rom = 8'b00011000;    // 5    **
            11'd390:    rom = 8'b00011000;    // 6    **
            11'd391:    rom = 8'b00011000;    // 7    **
            11'd392:    rom = 8'b00011000;    // 8    **
            11'd393:    rom = 8'b00011000;    // 9    **
            11'd394:    rom = 8'b00011000;    // a    **
            11'd395:    rom = 8'b00011000;    // b    **
            11'd396:    rom = 8'b00000000;    // c
            11'd397:    rom = 8'b00000000;    // d
            11'd398:    rom = 8'b00000000;    // e
            11'd399:    rom = 8'b00000000;    // f
   // code x19         
            11'd400:    rom = 8'b00000000;    // 0
            11'd401:    rom = 8'b00000000;    // 1
            11'd402:    rom = 8'b00011000;    // 2    **
            11'd403:    rom = 8'b00011000;    // 3    **
            11'd404:    rom = 8'b00011000;    // 4    **
            11'd405:    rom = 8'b00011000;    // 5    **
            11'd406:    rom = 8'b00011000;    // 6    **
            11'd407:    rom = 8'b00011000;    // 7    **
            11'd408:    rom = 8'b00011000;    // 8    **
            11'd409:    rom = 8'b01111110;    // 9  ******
            11'd410:    rom = 8'b00111100;    // a   ****
            11'd411:    rom = 8'b00011000;    // b    **
            11'd412:    rom = 8'b00000000;    // c
            11'd413:    rom = 8'b00000000;    // d
            11'd414:    rom = 8'b00000000;    // e
            11'd415:    rom = 8'b00000000;    // f
   // code x1a         
            11'd416:    rom = 8'b00000000;    // 0
            11'd417:    rom = 8'b00000000;    // 1
            11'd418:    rom = 8'b00000000;    // 2
            11'd419:    rom = 8'b00000000;    // 3
            11'd420:    rom = 8'b00000000;    // 4
            11'd421:    rom = 8'b00011000;    // 5    **
            11'd422:    rom = 8'b00001100;    // 6     **
            11'd423:    rom = 8'b11111110;    // 7 *******
            11'd424:    rom = 8'b00001100;    // 8     **
            11'd425:    rom = 8'b00011000;    // 9    **
            11'd426:    rom = 8'b00000000;    // a
            11'd427:    rom = 8'b00000000;    // b
            11'd428:    rom = 8'b00000000;    // c
            11'd429:    rom = 8'b00000000;    // d
            11'd430:    rom = 8'b00000000;    // e
            11'd431:    rom = 8'b00000000;    // f
   // code x1b         
            11'd432:    rom = 8'b00000000;    // 0
            11'd433:    rom = 8'b00000000;    // 1
            11'd434:    rom = 8'b00000000;    // 2
            11'd435:    rom = 8'b00000000;    // 3
            11'd436:    rom = 8'b00000000;    // 4
            11'd437:    rom = 8'b00110000;    // 5   **
            11'd438:    rom = 8'b01100000;    // 6  **
            11'd439:    rom = 8'b11111110;    // 7 *******
            11'd440:    rom = 8'b01100000;    // 8  **
            11'd441:    rom = 8'b00110000;    // 9   **
            11'd442:    rom = 8'b00000000;    // a
            11'd443:    rom = 8'b00000000;    // b
            11'd444:    rom = 8'b00000000;    // c
            11'd445:    rom = 8'b00000000;    // d
            11'd446:    rom = 8'b00000000;    // e
            11'd447:    rom = 8'b00000000;    // f
   // code x1c         
            11'd448:    rom = 8'b00000000;    // 0
            11'd449:    rom = 8'b00000000;    // 1
            11'd450:    rom = 8'b00000000;    // 2
            11'd451:    rom = 8'b00000000;    // 3
            11'd452:    rom = 8'b00000000;    // 4
            11'd453:    rom = 8'b00000000;    // 5
            11'd454:    rom = 8'b11000000;    // 6 **
            11'd455:    rom = 8'b11000000;    // 7 **
            11'd456:    rom = 8'b11000000;    // 8 **
            11'd457:    rom = 8'b11111110;    // 9 *******
            11'd458:    rom = 8'b00000000;    // a
            11'd459:    rom = 8'b00000000;    // b
            11'd460:    rom = 8'b00000000;    // c
            11'd461:    rom = 8'b00000000;    // d
            11'd462:    rom = 8'b00000000;    // e
            11'd463:    rom = 8'b00000000;    // f
   // code x1d         
            11'd464:    rom = 8'b00000000;    // 0
            11'd465:    rom = 8'b00000000;    // 1
            11'd466:    rom = 8'b00000000;    // 2
            11'd467:    rom = 8'b00000000;    // 3
            11'd468:    rom = 8'b00000000;    // 4
            11'd469:    rom = 8'b00100100;    // 5   *  *
            11'd470:    rom = 8'b01100110;    // 6  **  **
            11'd471:    rom = 8'b11111111;    // 7 ********
            11'd472:    rom = 8'b01100110;    // 8  **  **
            11'd473:    rom = 8'b00100100;    // 9   *  *
            11'd474:    rom = 8'b00000000;    // a
            11'd475:    rom = 8'b00000000;    // b
            11'd476:    rom = 8'b00000000;    // c
            11'd477:    rom = 8'b00000000;    // d
            11'd478:    rom = 8'b00000000;    // e
            11'd479:    rom = 8'b00000000;    // f
   // code x1e         
            11'd480:    rom = 8'b00000000;    // 0
            11'd481:    rom = 8'b00000000;    // 1
            11'd482:    rom = 8'b00000000;    // 2
            11'd483:    rom = 8'b00000000;    // 3
            11'd484:    rom = 8'b00010000;    // 4    *
            11'd485:    rom = 8'b00111000;    // 5   ***
            11'd486:    rom = 8'b00111000;    // 6   ***
            11'd487:    rom = 8'b01111100;    // 7  *****
            11'd488:    rom = 8'b01111100;    // 8  *****
            11'd489:    rom = 8'b11111110;    // 9 *******
            11'd490:    rom = 8'b11111110;    // a *******
            11'd491:    rom = 8'b00000000;    // b
            11'd492:    rom = 8'b00000000;    // c
            11'd493:    rom = 8'b00000000;    // d
            11'd494:    rom = 8'b00000000;    // e
            11'd495:    rom = 8'b00000000;    // f
   // code x1f         
            11'd496:    rom = 8'b00000000;    // 0
            11'd497:    rom = 8'b00000000;    // 1
            11'd498:    rom = 8'b00000000;    // 2
            11'd499:    rom = 8'b00000000;    // 3
            11'd500:    rom = 8'b11111110;    // 4 *******
            11'd501:    rom = 8'b11111110;    // 5 *******
            11'd502:    rom = 8'b01111100;    // 6  *****
            11'd503:    rom = 8'b01111100;    // 7  *****
            11'd504:    rom = 8'b00111000;    // 8   ***
            11'd505:    rom = 8'b00111000;    // 9   ***
            11'd506:    rom = 8'b00010000;    // a    *
            11'd507:    rom = 8'b00000000;    // b
            11'd508:    rom = 8'b00000000;    // c
            11'd509:    rom = 8'b00000000;    // d
            11'd510:    rom = 8'b00000000;    // e
            11'd511:    rom = 8'b00000000;    // f
   // code x20         
            11'd512:    rom = 8'b00000000;    // 0
            11'd513:    rom = 8'b00000000;    // 1
            11'd514:    rom = 8'b00000000;    // 2
            11'd515:    rom = 8'b00000000;    // 3
            11'd516:    rom = 8'b00000000;    // 4
            11'd517:    rom = 8'b00000000;    // 5
            11'd518:    rom = 8'b00000000;    // 6
            11'd519:    rom = 8'b00000000;    // 7
            11'd520:    rom = 8'b00000000;    // 8
            11'd521:    rom = 8'b00000000;    // 9
            11'd522:    rom = 8'b00000000;    // a
            11'd523:    rom = 8'b00000000;    // b
            11'd524:    rom = 8'b00000000;    // c
            11'd525:    rom = 8'b00000000;    // d
            11'd526:    rom = 8'b00000000;    // e
            11'd527:    rom = 8'b00000000;    // f
   // code x21         
            11'd528:    rom = 8'b00000000;    // 0
            11'd529:    rom = 8'b00000000;    // 1
            11'd530:    rom = 8'b00011000;    // 2    **
            11'd531:    rom = 8'b00111100;    // 3   ****
            11'd532:    rom = 8'b00111100;    // 4   ****
            11'd533:    rom = 8'b00111100;    // 5   ****
            11'd534:    rom = 8'b00011000;    // 6    **
            11'd535:    rom = 8'b00011000;    // 7    **
            11'd536:    rom = 8'b00011000;    // 8    **
            11'd537:    rom = 8'b00000000;    // 9
            11'd538:    rom = 8'b00011000;    // a    **
            11'd539:    rom = 8'b00011000;    // b    **
            11'd540:    rom = 8'b00000000;    // c
            11'd541:    rom = 8'b00000000;    // d
            11'd542:    rom = 8'b00000000;    // e
            11'd543:    rom = 8'b00000000;    // f
   // code x22         
            11'd544:    rom = 8'b00000000;    // 0
            11'd545:    rom = 8'b01100110;    // 1  **  **
            11'd546:    rom = 8'b01100110;    // 2  **  **
            11'd547:    rom = 8'b01100110;    // 3  **  **
            11'd548:    rom = 8'b00100100;    // 4   *  *
            11'd549:    rom = 8'b00000000;    // 5
            11'd550:    rom = 8'b00000000;    // 6
            11'd551:    rom = 8'b00000000;    // 7
            11'd552:    rom = 8'b00000000;    // 8
            11'd553:    rom = 8'b00000000;    // 9
            11'd554:    rom = 8'b00000000;    // a
            11'd555:    rom = 8'b00000000;    // b
            11'd556:    rom = 8'b00000000;    // c
            11'd557:    rom = 8'b00000000;    // d
            11'd558:    rom = 8'b00000000;    // e
            11'd559:    rom = 8'b00000000;    // f
   // code x23         
            11'd560:    rom = 8'b00000000;    // 0
            11'd561:    rom = 8'b00000000;    // 1
            11'd562:    rom = 8'b00000000;    // 2
            11'd563:    rom = 8'b01101100;    // 3  ** **
            11'd564:    rom = 8'b01101100;    // 4  ** **
            11'd565:    rom = 8'b11111110;    // 5 *******
            11'd566:    rom = 8'b01101100;    // 6  ** **
            11'd567:    rom = 8'b01101100;    // 7  ** **
            11'd568:    rom = 8'b01101100;    // 8  ** **
            11'd569:    rom = 8'b11111110;    // 9 *******
            11'd570:    rom = 8'b01101100;    // a  ** **
            11'd571:    rom = 8'b01101100;    // b  ** **
            11'd572:    rom = 8'b00000000;    // c
            11'd573:    rom = 8'b00000000;    // d
            11'd574:    rom = 8'b00000000;    // e
            11'd575:    rom = 8'b00000000;    // f
   // code x24         
            11'd576:    rom = 8'b00011000;    // 0     **
            11'd577:    rom = 8'b00011000;    // 1     **
            11'd578:    rom = 8'b01111100;    // 2   *****
            11'd579:    rom = 8'b11000110;    // 3  **   **
            11'd580:    rom = 8'b11000010;    // 4  **    *
            11'd581:    rom = 8'b11000000;    // 5  **
            11'd582:    rom = 8'b01111100;    // 6   *****
            11'd583:    rom = 8'b00000110;    // 7       **
            11'd584:    rom = 8'b00000110;    // 8       **
            11'd585:    rom = 8'b10000110;    // 9  *    **
            11'd586:    rom = 8'b11000110;    // a  **   **
            11'd587:    rom = 8'b01111100;    // b   *****
            11'd588:    rom = 8'b00011000;    // c     **
            11'd589:    rom = 8'b00011000;    // d     **
            11'd590:    rom = 8'b00000000;    // e
            11'd591:    rom = 8'b00000000;    // f
   // code x25         
            11'd592:    rom = 8'b00000000;    // 0
            11'd593:    rom = 8'b00000000;    // 1
            11'd594:    rom = 8'b00000000;    // 2
            11'd595:    rom = 8'b00000000;    // 3
            11'd596:    rom = 8'b11000010;    // 4 **    *
            11'd597:    rom = 8'b11000110;    // 5 **   **
            11'd598:    rom = 8'b00001100;    // 6     **
            11'd599:    rom = 8'b00011000;    // 7    **
            11'd600:    rom = 8'b00110000;    // 8   **
            11'd601:    rom = 8'b01100000;    // 9  **
            11'd602:    rom = 8'b11000110;    // a **   **
            11'd603:    rom = 8'b10000110;    // b *    **
            11'd604:    rom = 8'b00000000;    // c
            11'd605:    rom = 8'b00000000;    // d
            11'd606:    rom = 8'b00000000;    // e
            11'd607:    rom = 8'b00000000;    // f
   // code x26         
            11'd608:    rom = 8'b00000000;    // 0
            11'd609:    rom = 8'b00000000;    // 1
            11'd610:    rom = 8'b00111000;    // 2   ***
            11'd611:    rom = 8'b01101100;    // 3  ** **
            11'd612:    rom = 8'b01101100;    // 4  ** **
            11'd613:    rom = 8'b00111000;    // 5   ***
            11'd614:    rom = 8'b01110110;    // 6  *** **
            11'd615:    rom = 8'b11011100;    // 7 ** ***
            11'd616:    rom = 8'b11001100;    // 8 **  **
            11'd617:    rom = 8'b11001100;    // 9 **  **
            11'd618:    rom = 8'b11001100;    // a **  **
            11'd619:    rom = 8'b01110110;    // b  *** **
            11'd620:    rom = 8'b00000000;    // c
            11'd621:    rom = 8'b00000000;    // d
            11'd622:    rom = 8'b00000000;    // e
            11'd623:    rom = 8'b00000000;    // f
   // code x27         
            11'd624:    rom = 8'b00000000;    // 0
            11'd625:    rom = 8'b00110000;    // 1   **
            11'd626:    rom = 8'b00110000;    // 2   **
            11'd627:    rom = 8'b00110000;    // 3   **
            11'd628:    rom = 8'b01100000;    // 4  **
            11'd629:    rom = 8'b00000000;    // 5
            11'd630:    rom = 8'b00000000;    // 6
            11'd631:    rom = 8'b00000000;    // 7
            11'd632:    rom = 8'b00000000;    // 8
            11'd633:    rom = 8'b00000000;    // 9
            11'd634:    rom = 8'b00000000;    // a
            11'd635:    rom = 8'b00000000;    // b
            11'd636:    rom = 8'b00000000;    // c
            11'd637:    rom = 8'b00000000;    // d
            11'd638:    rom = 8'b00000000;    // e
            11'd639:    rom = 8'b00000000;    // f
   // code x28         
            11'd640:    rom = 8'b00000000;    // 0
            11'd641:    rom = 8'b00000000;    // 1
            11'd642:    rom = 8'b00001100;    // 2     **
            11'd643:    rom = 8'b00011000;    // 3    **
            11'd644:    rom = 8'b00110000;    // 4   **
            11'd645:    rom = 8'b00110000;    // 5   **
            11'd646:    rom = 8'b00110000;    // 6   **
            11'd647:    rom = 8'b00110000;    // 7   **
            11'd648:    rom = 8'b00110000;    // 8   **
            11'd649:    rom = 8'b00110000;    // 9   **
            11'd650:    rom = 8'b00011000;    // a    **
            11'd651:    rom = 8'b00001100;    // b     **
            11'd652:    rom = 8'b00000000;    // c
            11'd653:    rom = 8'b00000000;    // d
            11'd654:    rom = 8'b00000000;    // e
            11'd655:    rom = 8'b00000000;    // f
   // code x29         
            11'd656:    rom = 8'b00000000;    // 0
            11'd657:    rom = 8'b00000000;    // 1
            11'd658:    rom = 8'b00110000;    // 2   **
            11'd659:    rom = 8'b00011000;    // 3    **
            11'd660:    rom = 8'b00001100;    // 4     **
            11'd661:    rom = 8'b00001100;    // 5     **
            11'd662:    rom = 8'b00001100;    // 6     **
            11'd663:    rom = 8'b00001100;    // 7     **
            11'd664:    rom = 8'b00001100;    // 8     **
            11'd665:    rom = 8'b00001100;    // 9     **
            11'd666:    rom = 8'b00011000;    // a    **
            11'd667:    rom = 8'b00110000;    // b   **
            11'd668:    rom = 8'b00000000;    // c
            11'd669:    rom = 8'b00000000;    // d
            11'd670:    rom = 8'b00000000;    // e
            11'd671:    rom = 8'b00000000;    // f
   // code x2a         
            11'd672:    rom = 8'b00000000;    // 0
            11'd673:    rom = 8'b00000000;    // 1
            11'd674:    rom = 8'b00000000;    // 2
            11'd675:    rom = 8'b00000000;    // 3
            11'd676:    rom = 8'b00000000;    // 4
            11'd677:    rom = 8'b01100110;    // 5  **  **
            11'd678:    rom = 8'b00111100;    // 6   ****
            11'd679:    rom = 8'b11111111;    // 7 ********
            11'd680:    rom = 8'b00111100;    // 8   ****
            11'd681:    rom = 8'b01100110;    // 9  **  **
            11'd682:    rom = 8'b00000000;    // a
            11'd683:    rom = 8'b00000000;    // b
            11'd684:    rom = 8'b00000000;    // c
            11'd685:    rom = 8'b00000000;    // d
            11'd686:    rom = 8'b00000000;    // e
            11'd687:    rom = 8'b00000000;    // f
   // code x2b         
            11'd688:    rom = 8'b00000000;    // 0
            11'd689:    rom = 8'b00000000;    // 1
            11'd690:    rom = 8'b00000000;    // 2
            11'd691:    rom = 8'b00000000;    // 3
            11'd692:    rom = 8'b00000000;    // 4
            11'd693:    rom = 8'b00011000;    // 5    **
            11'd694:    rom = 8'b00011000;    // 6    **
            11'd695:    rom = 8'b01111110;    // 7  ******
            11'd696:    rom = 8'b00011000;    // 8    **
            11'd697:    rom = 8'b00011000;    // 9    **
            11'd698:    rom = 8'b00000000;    // a
            11'd699:    rom = 8'b00000000;    // b
            11'd700:    rom = 8'b00000000;    // c
            11'd701:    rom = 8'b00000000;    // d
            11'd702:    rom = 8'b00000000;    // e
            11'd703:    rom = 8'b00000000;    // f
   // code x2c         
            11'd704:    rom = 8'b00000000;    // 0
            11'd705:    rom = 8'b00000000;    // 1
            11'd706:    rom = 8'b00000000;    // 2
            11'd707:    rom = 8'b00000000;    // 3
            11'd708:    rom = 8'b00000000;    // 4
            11'd709:    rom = 8'b00000000;    // 5
            11'd710:    rom = 8'b00000000;    // 6
            11'd711:    rom = 8'b00000000;    // 7
            11'd712:    rom = 8'b00000000;    // 8
            11'd713:    rom = 8'b00011000;    // 9    **
            11'd714:    rom = 8'b00011000;    // a    **
            11'd715:    rom = 8'b00011000;    // b    **
            11'd716:    rom = 8'b00110000;    // c   **
            11'd717:    rom = 8'b00000000;    // d
            11'd718:    rom = 8'b00000000;    // e
            11'd719:    rom = 8'b00000000;    // f
   // code x2d         
            11'd720:    rom = 8'b00000000;    // 0
            11'd721:    rom = 8'b00000000;    // 1
            11'd722:    rom = 8'b00000000;    // 2
            11'd723:    rom = 8'b00000000;    // 3
            11'd724:    rom = 8'b00000000;    // 4
            11'd725:    rom = 8'b00000000;    // 5
            11'd726:    rom = 8'b00000000;    // 6
            11'd727:    rom = 8'b01111110;    // 7  ******
            11'd728:    rom = 8'b00000000;    // 8
            11'd729:    rom = 8'b00000000;    // 9
            11'd730:    rom = 8'b00000000;    // a
            11'd731:    rom = 8'b00000000;    // b
            11'd732:    rom = 8'b00000000;    // c
            11'd733:    rom = 8'b00000000;    // d
            11'd734:    rom = 8'b00000000;    // e
            11'd735:    rom = 8'b00000000;    // f
   // code x2e         
            11'd736:    rom = 8'b00000000;    // 0
            11'd737:    rom = 8'b00000000;    // 1
            11'd738:    rom = 8'b00000000;    // 2
            11'd739:    rom = 8'b00000000;    // 3
            11'd740:    rom = 8'b00000000;    // 4
            11'd741:    rom = 8'b00000000;    // 5
            11'd742:    rom = 8'b00000000;    // 6
            11'd743:    rom = 8'b00000000;    // 7
            11'd744:    rom = 8'b00000000;    // 8
            11'd745:    rom = 8'b00000000;    // 9
            11'd746:    rom = 8'b00011000;    // a    **
            11'd747:    rom = 8'b00011000;    // b    **
            11'd748:    rom = 8'b00000000;    // c
            11'd749:    rom = 8'b00000000;    // d
            11'd750:    rom = 8'b00000000;    // e
            11'd751:    rom = 8'b00000000;    // f
   // code x2f         
            11'd752:    rom = 8'b00000000;    // 0
            11'd753:    rom = 8'b00000000;    // 1
            11'd754:    rom = 8'b00000000;    // 2
            11'd755:    rom = 8'b00000000;    // 3
            11'd756:    rom = 8'b00000010;    // 4       *
            11'd757:    rom = 8'b00000110;    // 5      **
            11'd758:    rom = 8'b00001100;    // 6     **
            11'd759:    rom = 8'b00011000;    // 7    **
            11'd760:    rom = 8'b00110000;    // 8   **
            11'd761:    rom = 8'b01100000;    // 9  **
            11'd762:    rom = 8'b11000000;    // a **
            11'd763:    rom = 8'b10000000;    // b *
            11'd764:    rom = 8'b00000000;    // c
            11'd765:    rom = 8'b00000000;    // d
            11'd766:    rom = 8'b00000000;    // e
            11'd767:    rom = 8'b00000000;    // f
   // code x30         
            11'd768:    rom = 8'b00000000;    // 0
            11'd769:    rom = 8'b00000000;    // 1
            11'd770:    rom = 8'b01111100;    // 2  *****
            11'd771:    rom = 8'b11000110;    // 3 **   **
            11'd772:    rom = 8'b11000110;    // 4 **   **
            11'd773:    rom = 8'b11001110;    // 5 **  ***
            11'd774:    rom = 8'b11011110;    // 6 ** ****
            11'd775:    rom = 8'b11110110;    // 7 **** **
            11'd776:    rom = 8'b11100110;    // 8 ***  **
            11'd777:    rom = 8'b11000110;    // 9 **   **
            11'd778:    rom = 8'b11000110;    // a **   **
            11'd779:    rom = 8'b01111100;    // b  *****
            11'd780:    rom = 8'b00000000;    // c
            11'd781:    rom = 8'b00000000;    // d
            11'd782:    rom = 8'b00000000;    // e
            11'd783:    rom = 8'b00000000;    // f
   // code x31         
            11'd784:    rom = 8'b00000000;    // 0
            11'd785:    rom = 8'b00000000;    // 1
            11'd786:    rom = 8'b00011000;    // 2
            11'd787:    rom = 8'b00111000;    // 3
            11'd788:    rom = 8'b01111000;    // 4    **
            11'd789:    rom = 8'b00011000;    // 5   ***
            11'd790:    rom = 8'b00011000;    // 6  ****
            11'd791:    rom = 8'b00011000;    // 7    **
            11'd792:    rom = 8'b00011000;    // 8    **
            11'd793:    rom = 8'b00011000;    // 9    **
            11'd794:    rom = 8'b00011000;    // a    **
            11'd795:    rom = 8'b01111110;    // b    **
            11'd796:    rom = 8'b00000000;    // c    **
            11'd797:    rom = 8'b00000000;    // d  ******
            11'd798:    rom = 8'b00000000;    // e
            11'd799:    rom = 8'b00000000;    // f
   // code x32         
            11'd800:    rom = 8'b00000000;    // 0
            11'd801:    rom = 8'b00000000;    // 1
            11'd802:    rom = 8'b01111100;    // 2  *****
            11'd803:    rom = 8'b11000110;    // 3 **   **
            11'd804:    rom = 8'b00000110;    // 4      **
            11'd805:    rom = 8'b00001100;    // 5     **
            11'd806:    rom = 8'b00011000;    // 6    **
            11'd807:    rom = 8'b00110000;    // 7   **
            11'd808:    rom = 8'b01100000;    // 8  **
            11'd809:    rom = 8'b11000000;    // 9 **
            11'd810:    rom = 8'b11000110;    // a **   **
            11'd811:    rom = 8'b11111110;    // b *******
            11'd812:    rom = 8'b00000000;    // c
            11'd813:    rom = 8'b00000000;    // d
            11'd814:    rom = 8'b00000000;    // e
            11'd815:    rom = 8'b00000000;    // f
   // code x33         
            11'd816:    rom = 8'b00000000;    // 0
            11'd817:    rom = 8'b00000000;    // 1
            11'd818:    rom = 8'b01111100;    // 2  *****
            11'd819:    rom = 8'b11000110;    // 3 **   **
            11'd820:    rom = 8'b00000110;    // 4      **
            11'd821:    rom = 8'b00000110;    // 5      **
            11'd822:    rom = 8'b00111100;    // 6   ****
            11'd823:    rom = 8'b00000110;    // 7      **
            11'd824:    rom = 8'b00000110;    // 8      **
            11'd825:    rom = 8'b00000110;    // 9      **
            11'd826:    rom = 8'b11000110;    // a **   **
            11'd827:    rom = 8'b01111100;    // b  *****
            11'd828:    rom = 8'b00000000;    // c
            11'd829:    rom = 8'b00000000;    // d
            11'd830:    rom = 8'b00000000;    // e
            11'd831:    rom = 8'b00000000;    // f
   // code x34         
            11'd832:    rom = 8'b00000000;    // 0
            11'd833:    rom = 8'b00000000;    // 1
            11'd834:    rom = 8'b00001100;    // 2     **
            11'd835:    rom = 8'b00011100;    // 3    ***
            11'd836:    rom = 8'b00111100;    // 4   ****
            11'd837:    rom = 8'b01101100;    // 5  ** **
            11'd838:    rom = 8'b11001100;    // 6 **  **
            11'd839:    rom = 8'b11111110;    // 7 *******
            11'd840:    rom = 8'b00001100;    // 8     **
            11'd841:    rom = 8'b00001100;    // 9     **
            11'd842:    rom = 8'b00001100;    // a     **
            11'd843:    rom = 8'b00011110;    // b    ****
            11'd844:    rom = 8'b00000000;    // c
            11'd845:    rom = 8'b00000000;    // d
            11'd846:    rom = 8'b00000000;    // e
            11'd847:    rom = 8'b00000000;    // f
   // code x35         
            11'd848:    rom = 8'b00000000;    // 0
            11'd849:    rom = 8'b00000000;    // 1
            11'd850:    rom = 8'b11111110;    // 2 *******
            11'd851:    rom = 8'b11000000;    // 3 **
            11'd852:    rom = 8'b11000000;    // 4 **
            11'd853:    rom = 8'b11000000;    // 5 **
            11'd854:    rom = 8'b11111100;    // 6 ******
            11'd855:    rom = 8'b00000110;    // 7      **
            11'd856:    rom = 8'b00000110;    // 8      **
            11'd857:    rom = 8'b00000110;    // 9      **
            11'd858:    rom = 8'b11000110;    // a **   **
            11'd859:    rom = 8'b01111100;    // b  *****
            11'd860:    rom = 8'b00000000;    // c
            11'd861:    rom = 8'b00000000;    // d
            11'd862:    rom = 8'b00000000;    // e
            11'd863:    rom = 8'b00000000;    // f
   // code x36         
            11'd864:    rom = 8'b00000000;    // 0
            11'd865:    rom = 8'b00000000;    // 1
            11'd866:    rom = 8'b00111000;    // 2   ***
            11'd867:    rom = 8'b01100000;    // 3  **
            11'd868:    rom = 8'b11000000;    // 4 **
            11'd869:    rom = 8'b11000000;    // 5 **
            11'd870:    rom = 8'b11111100;    // 6 ******
            11'd871:    rom = 8'b11000110;    // 7 **   **
            11'd872:    rom = 8'b11000110;    // 8 **   **
            11'd873:    rom = 8'b11000110;    // 9 **   **
            11'd874:    rom = 8'b11000110;    // a **   **
            11'd875:    rom = 8'b01111100;    // b  *****
            11'd876:    rom = 8'b00000000;    // c
            11'd877:    rom = 8'b00000000;    // d
            11'd878:    rom = 8'b00000000;    // e
            11'd879:    rom = 8'b00000000;    // f
   // code x37         
            11'd880:    rom = 8'b00000000;    // 0
            11'd881:    rom = 8'b00000000;    // 1
            11'd882:    rom = 8'b11111110;    // 2 *******
            11'd883:    rom = 8'b11000110;    // 3 **   **
            11'd884:    rom = 8'b00000110;    // 4      **
            11'd885:    rom = 8'b00000110;    // 5      **
            11'd886:    rom = 8'b00001100;    // 6     **
            11'd887:    rom = 8'b00011000;    // 7    **
            11'd888:    rom = 8'b00110000;    // 8   **
            11'd889:    rom = 8'b00110000;    // 9   **
            11'd890:    rom = 8'b00110000;    // a   **
            11'd891:    rom = 8'b00110000;    // b   **
            11'd892:    rom = 8'b00000000;    // c
            11'd893:    rom = 8'b00000000;    // d
            11'd894:    rom = 8'b00000000;    // e
            11'd895:    rom = 8'b00000000;    // f
   // code x38         
            11'd896:    rom = 8'b00000000;    // 0
            11'd897:    rom = 8'b00000000;    // 1
            11'd898:    rom = 8'b01111100;    // 2  *****
            11'd899:    rom = 8'b11000110;    // 3 **   **
            11'd900:    rom = 8'b11000110;    // 4 **   **
            11'd901:    rom = 8'b11000110;    // 5 **   **
            11'd902:    rom = 8'b01111100;    // 6  *****
            11'd903:    rom = 8'b11000110;    // 7 **   **
            11'd904:    rom = 8'b11000110;    // 8 **   **
            11'd905:    rom = 8'b11000110;    // 9 **   **
            11'd906:    rom = 8'b11000110;    // a **   **
            11'd907:    rom = 8'b01111100;    // b  *****
            11'd908:    rom = 8'b00000000;    // c
            11'd909:    rom = 8'b00000000;    // d
            11'd910:    rom = 8'b00000000;    // e
            11'd911:    rom = 8'b00000000;    // f
   // code x39         
            11'd912:    rom = 8'b00000000;    // 0
            11'd913:    rom = 8'b00000000;    // 1
            11'd914:    rom = 8'b01111100;    // 2  *****
            11'd915:    rom = 8'b11000110;    // 3 **   **
            11'd916:    rom = 8'b11000110;    // 4 **   **
            11'd917:    rom = 8'b11000110;    // 5 **   **
            11'd918:    rom = 8'b01111110;    // 6  ******
            11'd919:    rom = 8'b00000110;    // 7      **
            11'd920:    rom = 8'b00000110;    // 8      **
            11'd921:    rom = 8'b00000110;    // 9      **
            11'd922:    rom = 8'b00001100;    // a     **
            11'd923:    rom = 8'b01111000;    // b  ****
            11'd924:    rom = 8'b00000000;    // c
            11'd925:    rom = 8'b00000000;    // d
            11'd926:    rom = 8'b00000000;    // e
            11'd927:    rom = 8'b00000000;    // f
   // code x3a         
            11'd928:    rom = 8'b00000000;    // 0
            11'd929:    rom = 8'b00000000;    // 1
            11'd930:    rom = 8'b00000000;    // 2
            11'd931:    rom = 8'b00000000;    // 3
            11'd932:    rom = 8'b00011000;    // 4    **
            11'd933:    rom = 8'b00011000;    // 5    **
            11'd934:    rom = 8'b00000000;    // 6
            11'd935:    rom = 8'b00000000;    // 7
            11'd936:    rom = 8'b00000000;    // 8
            11'd937:    rom = 8'b00011000;    // 9    **
            11'd938:    rom = 8'b00011000;    // a    **
            11'd939:    rom = 8'b00000000;    // b
            11'd940:    rom = 8'b00000000;    // c
            11'd941:    rom = 8'b00000000;    // d
            11'd942:    rom = 8'b00000000;    // e
            11'd943:    rom = 8'b00000000;    // f
   // code x3b         
            11'd944:    rom = 8'b00000000;    // 0
            11'd945:    rom = 8'b00000000;    // 1
            11'd946:    rom = 8'b00000000;    // 2
            11'd947:    rom = 8'b00000000;    // 3
            11'd948:    rom = 8'b00011000;    // 4    **
            11'd949:    rom = 8'b00011000;    // 5    **
            11'd950:    rom = 8'b00000000;    // 6
            11'd951:    rom = 8'b00000000;    // 7
            11'd952:    rom = 8'b00000000;    // 8
            11'd953:    rom = 8'b00011000;    // 9    **
            11'd954:    rom = 8'b00011000;    // a    **
            11'd955:    rom = 8'b00110000;    // b   **
            11'd956:    rom = 8'b00000000;    // c
            11'd957:    rom = 8'b00000000;    // d
            11'd958:    rom = 8'b00000000;    // e
            11'd959:    rom = 8'b00000000;    // f
   // code x3c         
            11'd960:    rom = 8'b00000000;    // 0
            11'd961:    rom = 8'b00000000;    // 1
            11'd962:    rom = 8'b00000000;    // 2
            11'd963:    rom = 8'b00000110;    // 3      **
            11'd964:    rom = 8'b00001100;    // 4     **
            11'd965:    rom = 8'b00011000;    // 5    **
            11'd966:    rom = 8'b00110000;    // 6   **
            11'd967:    rom = 8'b01100000;    // 7  **
            11'd968:    rom = 8'b00110000;    // 8   **
            11'd969:    rom = 8'b00011000;    // 9    **
            11'd970:    rom = 8'b00001100;    // a     **
            11'd971:    rom = 8'b00000110;    // b      **
            11'd972:    rom = 8'b00000000;    // c
            11'd973:    rom = 8'b00000000;    // d
            11'd974:    rom = 8'b00000000;    // e
            11'd975:    rom = 8'b00000000;    // f
   // code x3d         
            11'd976:    rom = 8'b00000000;    // 0
            11'd977:    rom = 8'b00000000;    // 1
            11'd978:    rom = 8'b00000000;    // 2
            11'd979:    rom = 8'b00000000;    // 3
            11'd980:    rom = 8'b00000000;    // 4
            11'd981:    rom = 8'b01111110;    // 5  ******
            11'd982:    rom = 8'b00000000;    // 6
            11'd983:    rom = 8'b00000000;    // 7
            11'd984:    rom = 8'b01111110;    // 8  ******
            11'd985:    rom = 8'b00000000;    // 9
            11'd986:    rom = 8'b00000000;    // a
            11'd987:    rom = 8'b00000000;    // b
            11'd988:    rom = 8'b00000000;    // c
            11'd989:    rom = 8'b00000000;    // d
            11'd990:    rom = 8'b00000000;    // e
            11'd991:    rom = 8'b00000000;    // f
   // code x3e         
            11'd992:    rom = 8'b00000000;    // 0
            11'd993:    rom = 8'b00000000;    // 1
            11'd994:    rom = 8'b00000000;    // 2
            11'd995:    rom = 8'b01100000;    // 3  **
            11'd996:    rom = 8'b00110000;    // 4   **
            11'd997:    rom = 8'b00011000;    // 5    **
            11'd998:    rom = 8'b00001100;    // 6     **
            11'd999:    rom = 8'b00000110;    // 7      **
            11'd1000:   rom = 8'b00001100;    // 8     **
            11'd1001:   rom = 8'b00011000;    // 9    **
            11'd1002:   rom = 8'b00110000;    // a   **
            11'd1003:   rom = 8'b01100000;    // b  **
            11'd1004:   rom = 8'b00000000;    // c
            11'd1005:   rom = 8'b00000000;    // d
            11'd1006:   rom = 8'b00000000;    // e
            11'd1007:   rom = 8'b00000000;    // f
   // code x3f
            11'd1008:   rom = 8'b00000000;    // 0
            11'd1009:   rom = 8'b00000000;    // 1
            11'd1010:   rom = 8'b01111100;    // 2  *****
            11'd1011:   rom = 8'b11000110;    // 3 **   **
            11'd1012:   rom = 8'b11000110;    // 4 **   **
            11'd1013:   rom = 8'b00001100;    // 5     **
            11'd1014:   rom = 8'b00011000;    // 6    **
            11'd1015:   rom = 8'b00011000;    // 7    **
            11'd1016:   rom = 8'b00011000;    // 8    **
            11'd1017:   rom = 8'b00000000;    // 9
            11'd1018:   rom = 8'b00011000;    // a    **
            11'd1019:   rom = 8'b00011000;    // b    **
            11'd1020:   rom = 8'b00000000;    // c
            11'd1021:   rom = 8'b00000000;    // d
            11'd1022:   rom = 8'b00000000;    // e
            11'd1023:   rom = 8'b00000000;    // f
   // code x40
            11'd1024:   rom = 8'b00000000;    // 0
            11'd1025:   rom = 8'b00000000;    // 1
            11'd1026:   rom = 8'b01111100;    // 2  *****
            11'd1027:   rom = 8'b11000110;    // 3 **   **
            11'd1028:   rom = 8'b11000110;    // 4 **   **
            11'd1029:   rom = 8'b11000110;    // 5 **   **
            11'd1030:   rom = 8'b11011110;    // 6 ** ****
            11'd1031:   rom = 8'b11011110;    // 7 ** ****
            11'd1032:   rom = 8'b11011110;    // 8 ** ****
            11'd1033:   rom = 8'b11011100;    // 9 ** ***
            11'd1034:   rom = 8'b11000000;    // a **
            11'd1035:   rom = 8'b01111100;    // b  *****
            11'd1036:   rom = 8'b00000000;    // c
            11'd1037:   rom = 8'b00000000;    // d
            11'd1038:   rom = 8'b00000000;    // e
            11'd1039:   rom = 8'b00000000;    // f
   // code x41
            11'd1040:   rom = 8'b00000000;    // 0
            11'd1041:   rom = 8'b00000000;    // 1
            11'd1042:   rom = 8'b00010000;    // 2    *
            11'd1043:   rom = 8'b00111000;    // 3   ***
            11'd1044:   rom = 8'b01101100;    // 4  ** **
            11'd1045:   rom = 8'b11000110;    // 5 **   **
            11'd1046:   rom = 8'b11000110;    // 6 **   **
            11'd1047:   rom = 8'b11111110;    // 7 *******
            11'd1048:   rom = 8'b11000110;    // 8 **   **
            11'd1049:   rom = 8'b11000110;    // 9 **   **
            11'd1050:   rom = 8'b11000110;    // a **   **
            11'd1051:   rom = 8'b11000110;    // b **   **
            11'd1052:   rom = 8'b00000000;    // c
            11'd1053:   rom = 8'b00000000;    // d
            11'd1054:   rom = 8'b00000000;    // e
            11'd1055:   rom = 8'b00000000;    // f
   // code x42
            11'd1056:   rom = 8'b00000000;    // 0
            11'd1057:   rom = 8'b00000000;    // 1
            11'd1058:   rom = 8'b11111100;    // 2 ******
            11'd1059:   rom = 8'b01100110;    // 3  **  **
            11'd1060:   rom = 8'b01100110;    // 4  **  **
            11'd1061:   rom = 8'b01100110;    // 5  **  **
            11'd1062:   rom = 8'b01111100;    // 6  *****
            11'd1063:   rom = 8'b01100110;    // 7  **  **
            11'd1064:   rom = 8'b01100110;    // 8  **  **
            11'd1065:   rom = 8'b01100110;    // 9  **  **
            11'd1066:   rom = 8'b01100110;    // a  **  **
            11'd1067:   rom = 8'b11111100;    // b ******
            11'd1068:   rom = 8'b00000000;    // c
            11'd1069:   rom = 8'b00000000;    // d
            11'd1070:   rom = 8'b00000000;    // e
            11'd1071:   rom = 8'b00000000;    // f
   // code x43
            11'd1072:   rom = 8'b00000000;    // 0
            11'd1073:   rom = 8'b00000000;    // 1
            11'd1074:   rom = 8'b00111100;    // 2   ****
            11'd1075:   rom = 8'b01100110;    // 3  **  **
            11'd1076:   rom = 8'b11000010;    // 4 **    *
            11'd1077:   rom = 8'b11000000;    // 5 **
            11'd1078:   rom = 8'b11000000;    // 6 **
            11'd1079:   rom = 8'b11000000;    // 7 **
            11'd1080:   rom = 8'b11000000;    // 8 **
            11'd1081:   rom = 8'b11000010;    // 9 **    *
            11'd1082:   rom = 8'b01100110;    // a  **  **
            11'd1083:   rom = 8'b00111100;    // b   ****
            11'd1084:   rom = 8'b00000000;    // c
            11'd1085:   rom = 8'b00000000;    // d
            11'd1086:   rom = 8'b00000000;    // e
            11'd1087:   rom = 8'b00000000;    // f
   // code x44
            11'd1088:   rom = 8'b00000000;    // 0
            11'd1089:   rom = 8'b00000000;    // 1
            11'd1090:   rom = 8'b11111000;    // 2 *****
            11'd1091:   rom = 8'b01101100;    // 3  ** **
            11'd1092:   rom = 8'b01100110;    // 4  **  **
            11'd1093:   rom = 8'b01100110;    // 5  **  **
            11'd1094:   rom = 8'b01100110;    // 6  **  **
            11'd1095:   rom = 8'b01100110;    // 7  **  **
            11'd1096:   rom = 8'b01100110;    // 8  **  **
            11'd1097:   rom = 8'b01100110;    // 9  **  **
            11'd1098:   rom = 8'b01101100;    // a  ** **
            11'd1099:   rom = 8'b11111000;    // b *****
            11'd1100:   rom = 8'b00000000;    // c
            11'd1101:   rom = 8'b00000000;    // d
            11'd1102:   rom = 8'b00000000;    // e
            11'd1103:   rom = 8'b00000000;    // f
   // code x45
            11'd1104:   rom = 8'b00000000;    // 0
            11'd1105:   rom = 8'b00000000;    // 1
            11'd1106:   rom = 8'b11111110;    // 2 *******
            11'd1107:   rom = 8'b01100110;    // 3  **  **
            11'd1108:   rom = 8'b01100010;    // 4  **   *
            11'd1109:   rom = 8'b01101000;    // 5  ** *
            11'd1110:   rom = 8'b01111000;    // 6  ****
            11'd1111:   rom = 8'b01101000;    // 7  ** *
            11'd1112:   rom = 8'b01100000;    // 8  **
            11'd1113:   rom = 8'b01100010;    // 9  **   *
            11'd1114:   rom = 8'b01100110;    // a  **  **
            11'd1115:   rom = 8'b11111110;    // b *******
            11'd1116:   rom = 8'b00000000;    // c
            11'd1117:   rom = 8'b00000000;    // d
            11'd1118:   rom = 8'b00000000;    // e
            11'd1119:   rom = 8'b00000000;    // f
   // code x46
            11'd1120:   rom = 8'b00000000;    // 0
            11'd1121:   rom = 8'b00000000;    // 1
            11'd1122:   rom = 8'b11111110;    // 2 *******
            11'd1123:   rom = 8'b01100110;    // 3  **  **
            11'd1124:   rom = 8'b01100010;    // 4  **   *
            11'd1125:   rom = 8'b01101000;    // 5  ** *
            11'd1126:   rom = 8'b01111000;    // 6  ****
            11'd1127:   rom = 8'b01101000;    // 7  ** *
            11'd1128:   rom = 8'b01100000;    // 8  **
            11'd1129:   rom = 8'b01100000;    // 9  **
            11'd1130:   rom = 8'b01100000;    // a  **
            11'd1131:   rom = 8'b11110000;    // b ****
            11'd1132:   rom = 8'b00000000;    // c
            11'd1133:   rom = 8'b00000000;    // d
            11'd1134:   rom = 8'b00000000;    // e
            11'd1135:   rom = 8'b00000000;    // f
   // code x47
            11'd1136:   rom = 8'b00000000;    // 0
            11'd1137:   rom = 8'b00000000;    // 1
            11'd1138:   rom = 8'b00111100;    // 2   ****
            11'd1139:   rom = 8'b01100110;    // 3  **  **
            11'd1140:   rom = 8'b11000010;    // 4 **    *
            11'd1141:   rom = 8'b11000000;    // 5 **
            11'd1142:   rom = 8'b11000000;    // 6 **
            11'd1143:   rom = 8'b11011110;    // 7 ** ****
            11'd1144:   rom = 8'b11000110;    // 8 **   **
            11'd1145:   rom = 8'b11000110;    // 9 **   **
            11'd1146:   rom = 8'b01100110;    // a  **  **
            11'd1147:   rom = 8'b00111010;    // b   *** *
            11'd1148:   rom = 8'b00000000;    // c
            11'd1149:   rom = 8'b00000000;    // d
            11'd1150:   rom = 8'b00000000;    // e
            11'd1151:   rom = 8'b00000000;    // f
   // code x48
            11'd1152:   rom = 8'b00000000;    // 0
            11'd1153:   rom = 8'b00000000;    // 1
            11'd1154:   rom = 8'b11000110;    // 2 **   **
            11'd1155:   rom = 8'b11000110;    // 3 **   **
            11'd1156:   rom = 8'b11000110;    // 4 **   **
            11'd1157:   rom = 8'b11000110;    // 5 **   **
            11'd1158:   rom = 8'b11111110;    // 6 *******
            11'd1159:   rom = 8'b11000110;    // 7 **   **
            11'd1160:   rom = 8'b11000110;    // 8 **   **
            11'd1161:   rom = 8'b11000110;    // 9 **   **
            11'd1162:   rom = 8'b11000110;    // a **   **
            11'd1163:   rom = 8'b11000110;    // b **   **
            11'd1164:   rom = 8'b00000000;    // c
            11'd1165:   rom = 8'b00000000;    // d
            11'd1166:   rom = 8'b00000000;    // e
            11'd1167:   rom = 8'b00000000;    // f
   // code x49
            11'd1168:   rom = 8'b00000000;    // 0
            11'd1169:   rom = 8'b00000000;    // 1
            11'd1170:   rom = 8'b00111100;    // 2   ****
            11'd1171:   rom = 8'b00011000;    // 3    **
            11'd1172:   rom = 8'b00011000;    // 4    **
            11'd1173:   rom = 8'b00011000;    // 5    **
            11'd1174:   rom = 8'b00011000;    // 6    **
            11'd1175:   rom = 8'b00011000;    // 7    **
            11'd1176:   rom = 8'b00011000;    // 8    **
            11'd1177:   rom = 8'b00011000;    // 9    **
            11'd1178:   rom = 8'b00011000;    // a    **
            11'd1179:   rom = 8'b00111100;    // b   ****
            11'd1180:   rom = 8'b00000000;    // c
            11'd1181:   rom = 8'b00000000;    // d
            11'd1182:   rom = 8'b00000000;    // e
            11'd1183:   rom = 8'b00000000;    // f
   // code x4a
            11'd1184:   rom = 8'b00000000;    // 0
            11'd1185:   rom = 8'b00000000;    // 1
            11'd1186:   rom = 8'b00011110;    // 2    ****
            11'd1187:   rom = 8'b00001100;    // 3     **
            11'd1188:   rom = 8'b00001100;    // 4     **
            11'd1189:   rom = 8'b00001100;    // 5     **
            11'd1190:   rom = 8'b00001100;    // 6     **
            11'd1191:   rom = 8'b00001100;    // 7     **
            11'd1192:   rom = 8'b11001100;    // 8 **  **
            11'd1193:   rom = 8'b11001100;    // 9 **  **
            11'd1194:   rom = 8'b11001100;    // a **  **
            11'd1195:   rom = 8'b01111000;    // b  ****
            11'd1196:   rom = 8'b00000000;    // c
            11'd1197:   rom = 8'b00000000;    // d
            11'd1198:   rom = 8'b00000000;    // e
            11'd1199:   rom = 8'b00000000;    // f
   // code x4b
            11'd1200:   rom = 8'b00000000;    // 0
            11'd1201:   rom = 8'b00000000;    // 1
            11'd1202:   rom = 8'b11100110;    // 2 ***  **
            11'd1203:   rom = 8'b01100110;    // 3  **  **
            11'd1204:   rom = 8'b01100110;    // 4  **  **
            11'd1205:   rom = 8'b01101100;    // 5  ** **
            11'd1206:   rom = 8'b01111000;    // 6  ****
            11'd1207:   rom = 8'b01111000;    // 7  ****
            11'd1208:   rom = 8'b01101100;    // 8  ** **
            11'd1209:   rom = 8'b01100110;    // 9  **  **
            11'd1210:   rom = 8'b01100110;    // a  **  **
            11'd1211:   rom = 8'b11100110;    // b ***  **
            11'd1212:   rom = 8'b00000000;    // c
            11'd1213:   rom = 8'b00000000;    // d
            11'd1214:   rom = 8'b00000000;    // e
            11'd1215:   rom = 8'b00000000;    // f
   // code x4c
            11'd1216:   rom = 8'b00000000;    // 0
            11'd1217:   rom = 8'b00000000;    // 1
            11'd1218:   rom = 8'b11110000;    // 2 ****
            11'd1219:   rom = 8'b01100000;    // 3  **
            11'd1220:   rom = 8'b01100000;    // 4  **
            11'd1221:   rom = 8'b01100000;    // 5  **
            11'd1222:   rom = 8'b01100000;    // 6  **
            11'd1223:   rom = 8'b01100000;    // 7  **
            11'd1224:   rom = 8'b01100000;    // 8  **
            11'd1225:   rom = 8'b01100010;    // 9  **   *
            11'd1226:   rom = 8'b01100110;    // a  **  **
            11'd1227:   rom = 8'b11111110;    // b *******
            11'd1228:   rom = 8'b00000000;    // c
            11'd1229:   rom = 8'b00000000;    // d
            11'd1230:   rom = 8'b00000000;    // e
            11'd1231:   rom = 8'b00000000;    // f
   // code x4d
            11'd1232:   rom = 8'b00000000;    // 0
            11'd1233:   rom = 8'b00000000;    // 1
            11'd1234:   rom = 8'b11000011;    // 2 **    **
            11'd1235:   rom = 8'b11100111;    // 3 ***  ***
            11'd1236:   rom = 8'b11111111;    // 4 ********
            11'd1237:   rom = 8'b11111111;    // 5 ********
            11'd1238:   rom = 8'b11011011;    // 6 ** ** **
            11'd1239:   rom = 8'b11000011;    // 7 **    **
            11'd1240:   rom = 8'b11000011;    // 8 **    **
            11'd1241:   rom = 8'b11000011;    // 9 **    **
            11'd1242:   rom = 8'b11000011;    // a **    **
            11'd1243:   rom = 8'b11000011;    // b **    **
            11'd1244:   rom = 8'b00000000;    // c
            11'd1245:   rom = 8'b00000000;    // d
            11'd1246:   rom = 8'b00000000;    // e
            11'd1247:   rom = 8'b00000000;    // f
   // code x4e
            11'd1248:   rom = 8'b00000000;    // 0
            11'd1249:   rom = 8'b00000000;    // 1
            11'd1250:   rom = 8'b11000110;    // 2 **   **
            11'd1251:   rom = 8'b11100110;    // 3 ***  **
            11'd1252:   rom = 8'b11110110;    // 4 **** **
            11'd1253:   rom = 8'b11111110;    // 5 *******
            11'd1254:   rom = 8'b11011110;    // 6 ** ****
            11'd1255:   rom = 8'b11001110;    // 7 **  ***
            11'd1256:   rom = 8'b11000110;    // 8 **   **
            11'd1257:   rom = 8'b11000110;    // 9 **   **
            11'd1258:   rom = 8'b11000110;    // a **   **
            11'd1259:   rom = 8'b11000110;    // b **   **
            11'd1260:   rom = 8'b00000000;    // c
            11'd1261:   rom = 8'b00000000;    // d
            11'd1262:   rom = 8'b00000000;    // e
            11'd1263:   rom = 8'b00000000;    // f
   // code x4f
            11'd1264:   rom = 8'b00000000;    // 0
            11'd1265:   rom = 8'b00000000;    // 1
            11'd1266:   rom = 8'b01111100;    // 2  *****
            11'd1267:   rom = 8'b11000110;    // 3 **   **
            11'd1268:   rom = 8'b11000110;    // 4 **   **
            11'd1269:   rom = 8'b11000110;    // 5 **   **
            11'd1270:   rom = 8'b11000110;    // 6 **   **
            11'd1271:   rom = 8'b11000110;    // 7 **   **
            11'd1272:   rom = 8'b11000110;    // 8 **   **
            11'd1273:   rom = 8'b11000110;    // 9 **   **
            11'd1274:   rom = 8'b11000110;    // a **   **
            11'd1275:   rom = 8'b01111100;    // b  *****
            11'd1276:   rom = 8'b00000000;    // c
            11'd1277:   rom = 8'b00000000;    // d
            11'd1278:   rom = 8'b00000000;    // e
            11'd1279:   rom = 8'b00000000;    // f
   // code x50
            11'd1280:   rom = 8'b00000000;    // 0
            11'd1281:   rom = 8'b00000000;    // 1
            11'd1282:   rom = 8'b11111100;    // 2 ******
            11'd1283:   rom = 8'b01100110;    // 3  **  **
            11'd1284:   rom = 8'b01100110;    // 4  **  **
            11'd1285:   rom = 8'b01100110;    // 5  **  **
            11'd1286:   rom = 8'b01111100;    // 6  *****
            11'd1287:   rom = 8'b01100000;    // 7  **
            11'd1288:   rom = 8'b01100000;    // 8  **
            11'd1289:   rom = 8'b01100000;    // 9  **
            11'd1290:   rom = 8'b01100000;    // a  **
            11'd1291:   rom = 8'b11110000;    // b ****
            11'd1292:   rom = 8'b00000000;    // c
            11'd1293:   rom = 8'b00000000;    // d
            11'd1294:   rom = 8'b00000000;    // e
            11'd1295:   rom = 8'b00000000;    // f
   // code x510
            11'd1296:   rom = 8'b00000000;    // 0
            11'd1297:   rom = 8'b00000000;    // 1
            11'd1298:   rom = 8'b01111100;    // 2  *****
            11'd1299:   rom = 8'b11000110;    // 3 **   **
            11'd1300:   rom = 8'b11000110;    // 4 **   **
            11'd1301:   rom = 8'b11000110;    // 5 **   **
            11'd1302:   rom = 8'b11000110;    // 6 **   **
            11'd1303:   rom = 8'b11000110;    // 7 **   **
            11'd1304:   rom = 8'b11000110;    // 8 **   **
            11'd1305:   rom = 8'b11010110;    // 9 ** * **
            11'd1306:   rom = 8'b11011110;    // a ** ****
            11'd1307:   rom = 8'b01111100;    // b  *****
            11'd1308:   rom = 8'b00001100;    // c     **
            11'd1309:   rom = 8'b00001110;    // d     ***
            11'd1310:   rom = 8'b00000000;    // e
            11'd1311:   rom = 8'b00000000;    // f
   // code x52
            11'd1312:   rom = 8'b00000000;    // 0
            11'd1313:   rom = 8'b00000000;    // 1
            11'd1314:   rom = 8'b11111100;    // 2 ******
            11'd1315:   rom = 8'b01100110;    // 3  **  **
            11'd1316:   rom = 8'b01100110;    // 4  **  **
            11'd1317:   rom = 8'b01100110;    // 5  **  **
            11'd1318:   rom = 8'b01111100;    // 6  *****
            11'd1319:   rom = 8'b01101100;    // 7  ** **
            11'd1320:   rom = 8'b01100110;    // 8  **  **
            11'd1321:   rom = 8'b01100110;    // 9  **  **
            11'd1322:   rom = 8'b01100110;    // a  **  **
            11'd1323:   rom = 8'b11100110;    // b ***  **
            11'd1324:   rom = 8'b00000000;    // c
            11'd1325:   rom = 8'b00000000;    // d
            11'd1326:   rom = 8'b00000000;    // e
            11'd1327:   rom = 8'b00000000;    // f
   // code x53
            11'd1328:   rom = 8'b00000000;    // 0
            11'd1329:   rom = 8'b00000000;    // 1
            11'd1330:   rom = 8'b01111100;    // 2  *****
            11'd1331:   rom = 8'b11000110;    // 3 **   **
            11'd1332:   rom = 8'b11000110;    // 4 **   **
            11'd1333:   rom = 8'b01100000;    // 5  **
            11'd1334:   rom = 8'b00111000;    // 6   ***
            11'd1335:   rom = 8'b00001100;    // 7     **
            11'd1336:   rom = 8'b00000110;    // 8      **
            11'd1337:   rom = 8'b11000110;    // 9 **   **
            11'd1338:   rom = 8'b11000110;    // a **   **
            11'd1339:   rom = 8'b01111100;    // b  *****
            11'd1340:   rom = 8'b00000000;    // c
            11'd1341:   rom = 8'b00000000;    // d
            11'd1342:   rom = 8'b00000000;    // e
            11'd1343:   rom = 8'b00000000;    // f
   // code x54
            11'd1344:   rom = 8'b00000000;    // 0
            11'd1345:   rom = 8'b00000000;    // 1
            11'd1346:   rom = 8'b11111111;    // 2 ********
            11'd1347:   rom = 8'b11011011;    // 3 ** ** **
            11'd1348:   rom = 8'b10011001;    // 4 *  **  *
            11'd1349:   rom = 8'b00011000;    // 5    **
            11'd1350:   rom = 8'b00011000;    // 6    **
            11'd1351:   rom = 8'b00011000;    // 7    **
            11'd1352:   rom = 8'b00011000;    // 8    **
            11'd1353:   rom = 8'b00011000;    // 9    **
            11'd1354:   rom = 8'b00011000;    // a    **
            11'd1355:   rom = 8'b00111100;    // b   ****
            11'd1356:   rom = 8'b00000000;    // c
            11'd1357:   rom = 8'b00000000;    // d
            11'd1358:   rom = 8'b00000000;    // e
            11'd1359:   rom = 8'b00000000;    // f
   // code x55
            11'd1360:   rom = 8'b00000000;    // 0
            11'd1361:   rom = 8'b00000000;    // 1
            11'd1362:   rom = 8'b11000110;    // 2 **   **
            11'd1363:   rom = 8'b11000110;    // 3 **   **
            11'd1364:   rom = 8'b11000110;    // 4 **   **
            11'd1365:   rom = 8'b11000110;    // 5 **   **
            11'd1366:   rom = 8'b11000110;    // 6 **   **
            11'd1367:   rom = 8'b11000110;    // 7 **   **
            11'd1368:   rom = 8'b11000110;    // 8 **   **
            11'd1369:   rom = 8'b11000110;    // 9 **   **
            11'd1370:   rom = 8'b11000110;    // a **   **
            11'd1371:   rom = 8'b01111100;    // b  *****
            11'd1372:   rom = 8'b00000000;    // c
            11'd1373:   rom = 8'b00000000;    // d
            11'd1374:   rom = 8'b00000000;    // e
            11'd1375:   rom = 8'b00000000;    // f
   // code x56
            11'd1376:   rom = 8'b00000000;    // 0
            11'd1377:   rom = 8'b00000000;    // 1
            11'd1378:   rom = 8'b11000011;    // 2 **    **
            11'd1379:   rom = 8'b11000011;    // 3 **    **
            11'd1380:   rom = 8'b11000011;    // 4 **    **
            11'd1381:   rom = 8'b11000011;    // 5 **    **
            11'd1382:   rom = 8'b11000011;    // 6 **    **
            11'd1383:   rom = 8'b11000011;    // 7 **    **
            11'd1384:   rom = 8'b11000011;    // 8 **    **
            11'd1385:   rom = 8'b01100110;    // 9  **  **
            11'd1386:   rom = 8'b00111100;    // a   ****
            11'd1387:   rom = 8'b00011000;    // b    **
            11'd1388:   rom = 8'b00000000;    // c
            11'd1389:   rom = 8'b00000000;    // d
            11'd1390:   rom = 8'b00000000;    // e
            11'd1391:   rom = 8'b00000000;    // f
   // code x57
            11'd1392:   rom = 8'b00000000;    // 0
            11'd1393:   rom = 8'b00000000;    // 1
            11'd1394:   rom = 8'b11000011;    // 2 **    **
            11'd1395:   rom = 8'b11000011;    // 3 **    **
            11'd1396:   rom = 8'b11000011;    // 4 **    **
            11'd1397:   rom = 8'b11000011;    // 5 **    **
            11'd1398:   rom = 8'b11000011;    // 6 **    **
            11'd1399:   rom = 8'b11011011;    // 7 ** ** **
            11'd1400:   rom = 8'b11011011;    // 8 ** ** **
            11'd1401:   rom = 8'b11111111;    // 9 ********
            11'd1402:   rom = 8'b01100110;    // a  **  **
            11'd1403:   rom = 8'b01100110;    // b  **  **
            11'd1404:   rom = 8'b00000000;    // c
            11'd1405:   rom = 8'b00000000;    // d
            11'd1406:   rom = 8'b00000000;    // e
            11'd1407:   rom = 8'b00000000;    // f

   // code x58
            11'd1408:   rom = 8'b00000000;    // 0
            11'd1409:   rom = 8'b00000000;    // 1
            11'd1410:   rom = 8'b11000011;    // 2 **    **
            11'd1411:   rom = 8'b11000011;    // 3 **    **
            11'd1412:   rom = 8'b01100110;    // 4  **  **
            11'd1413:   rom = 8'b00111100;    // 5   ****
            11'd1414:   rom = 8'b00011000;    // 6    **
            11'd1415:   rom = 8'b00011000;    // 7    **
            11'd1416:   rom = 8'b00111100;    // 8   ****
            11'd1417:   rom = 8'b01100110;    // 9  **  **
            11'd1418:   rom = 8'b11000011;    // a **    **
            11'd1419:   rom = 8'b11000011;    // b **    **
            11'd1420:   rom = 8'b00000000;    // c
            11'd1421:   rom = 8'b00000000;    // d
            11'd1422:   rom = 8'b00000000;    // e
            11'd1423:   rom = 8'b00000000;    // f
   // code x59
            11'd1424:   rom = 8'b00000000;    // 0
            11'd1425:   rom = 8'b00000000;    // 1
            11'd1426:   rom = 8'b11000011;    // 2 **    **
            11'd1427:   rom = 8'b11000011;    // 3 **    **
            11'd1428:   rom = 8'b11000011;    // 4 **    **
            11'd1429:   rom = 8'b01100110;    // 5  **  **
            11'd1430:   rom = 8'b00111100;    // 6   ****
            11'd1431:   rom = 8'b00011000;    // 7    **
            11'd1432:   rom = 8'b00011000;    // 8    **
            11'd1433:   rom = 8'b00011000;    // 9    **
            11'd1434:   rom = 8'b00011000;    // a    **
            11'd1435:   rom = 8'b00111100;    // b   ****
            11'd1436:   rom = 8'b00000000;    // c
            11'd1437:   rom = 8'b00000000;    // d
            11'd1438:   rom = 8'b00000000;    // e
            11'd1439:   rom = 8'b00000000;    // f
   // code x5a
            11'd1440:   rom = 8'b00000000;    // 0
            11'd1441:   rom = 8'b00000000;    // 1
            11'd1442:   rom = 8'b11111111;    // 2 ********
            11'd1443:   rom = 8'b11000011;    // 3 **    **
            11'd1444:   rom = 8'b10000110;    // 4 *    **
            11'd1445:   rom = 8'b00001100;    // 5     **
            11'd1446:   rom = 8'b00011000;    // 6    **
            11'd1447:   rom = 8'b00110000;    // 7   **
            11'd1448:   rom = 8'b01100000;    // 8  **
            11'd1449:   rom = 8'b11000001;    // 9 **     *
            11'd1450:   rom = 8'b11000011;    // a **    **
            11'd1451:   rom = 8'b11111111;    // b ********
            11'd1452:   rom = 8'b00000000;    // c
            11'd1453:   rom = 8'b00000000;    // d
            11'd1454:   rom = 8'b00000000;    // e
            11'd1455:   rom = 8'b00000000;    // f
   // code x5b
            11'd1456:   rom = 8'b00000000;    // 0
            11'd1457:   rom = 8'b00000000;    // 1
            11'd1458:   rom = 8'b00111100;    // 2   ****
            11'd1459:   rom = 8'b00110000;    // 3   **
            11'd1460:   rom = 8'b00110000;    // 4   **
            11'd1461:   rom = 8'b00110000;    // 5   **
            11'd1462:   rom = 8'b00110000;    // 6   **
            11'd1463:   rom = 8'b00110000;    // 7   **
            11'd1464:   rom = 8'b00110000;    // 8   **
            11'd1465:   rom = 8'b00110000;    // 9   **
            11'd1466:   rom = 8'b00110000;    // a   **
            11'd1467:   rom = 8'b00111100;    // b   ****
            11'd1468:   rom = 8'b00000000;    // c
            11'd1469:   rom = 8'b00000000;    // d
            11'd1470:   rom = 8'b00000000;    // e
            11'd1471:   rom = 8'b00000000;    // f
   // code x5c
            11'd1472:   rom = 8'b00000000;    // 0
            11'd1473:   rom = 8'b00000000;    // 1
            11'd1474:   rom = 8'b00000000;    // 2
            11'd1475:   rom = 8'b10000000;    // 3 *
            11'd1476:   rom = 8'b11000000;    // 4 **
            11'd1477:   rom = 8'b11100000;    // 5 ***
            11'd1478:   rom = 8'b01110000;    // 6  ***
            11'd1479:   rom = 8'b00111000;    // 7   ***
            11'd1480:   rom = 8'b00011100;    // 8    ***
            11'd1481:   rom = 8'b00001110;    // 9     ***
            11'd1482:   rom = 8'b00000110;    // a      **
            11'd1483:   rom = 8'b00000010;    // b       *
            11'd1484:   rom = 8'b00000000;    // c
            11'd1485:   rom = 8'b00000000;    // d
            11'd1486:   rom = 8'b00000000;    // e
            11'd1487:   rom = 8'b00000000;    // f
   // code x5d
            11'd1488:   rom = 8'b00000000;    // 0
            11'd1489:   rom = 8'b00000000;    // 1
            11'd1490:   rom = 8'b00111100;    // 2   ****
            11'd1491:   rom = 8'b00001100;    // 3     **
            11'd1492:   rom = 8'b00001100;    // 4     **
            11'd1493:   rom = 8'b00001100;    // 5     **
            11'd1494:   rom = 8'b00001100;    // 6     **
            11'd1495:   rom = 8'b00001100;    // 7     **
            11'd1496:   rom = 8'b00001100;    // 8     **
            11'd1497:   rom = 8'b00001100;    // 9     **
            11'd1498:   rom = 8'b00001100;    // a     **
            11'd1499:   rom = 8'b00111100;    // b   ****
            11'd1500:   rom = 8'b00000000;    // c
            11'd1501:   rom = 8'b00000000;    // d
            11'd1502:   rom = 8'b00000000;    // e
            11'd1503:   rom = 8'b00000000;    // f
   // code x5e
            11'd1504:   rom = 8'b00010000;    // 0    *
            11'd1505:   rom = 8'b00111000;    // 1   ***
            11'd1506:   rom = 8'b01101100;    // 2  ** **
            11'd1507:   rom = 8'b11000110;    // 3 **   **
            11'd1508:   rom = 8'b00000000;    // 4
            11'd1509:   rom = 8'b00000000;    // 5
            11'd1510:   rom = 8'b00000000;    // 6
            11'd1511:   rom = 8'b00000000;    // 7
            11'd1512:   rom = 8'b00000000;    // 8
            11'd1513:   rom = 8'b00000000;    // 9
            11'd1514:   rom = 8'b00000000;    // a
            11'd1515:   rom = 8'b00000000;    // b
            11'd1516:   rom = 8'b00000000;    // c
            11'd1517:   rom = 8'b00000000;    // d
            11'd1518:   rom = 8'b00000000;    // e
            11'd1519:   rom = 8'b00000000;    // f
   // code x5f
            11'd1520:   rom = 8'b00000000;    // 0
            11'd1521:   rom = 8'b00000000;    // 1
            11'd1522:   rom = 8'b00000000;    // 2
            11'd1523:   rom = 8'b00000000;    // 3
            11'd1524:   rom = 8'b00000000;    // 4
            11'd1525:   rom = 8'b00000000;    // 5
            11'd1526:   rom = 8'b00000000;    // 6
            11'd1527:   rom = 8'b00000000;    // 7
            11'd1528:   rom = 8'b00000000;    // 8
            11'd1529:   rom = 8'b00000000;    // 9
            11'd1530:   rom = 8'b00000000;    // a
            11'd1531:   rom = 8'b00000000;    // b
            11'd1532:   rom = 8'b00000000;    // c
            11'd1533:   rom = 8'b11111111;    // d ********
            11'd1534:   rom = 8'b00000000;    // e
            11'd1535:   rom = 8'b00000000;    // f
   // code x60
            11'd1536:   rom = 8'b00110000;    // 0   **
            11'd1537:   rom = 8'b00110000;    // 1   **
            11'd1538:   rom = 8'b00011000;    // 2    **
            11'd1539:   rom = 8'b00000000;    // 3
            11'd1540:   rom = 8'b00000000;    // 4
            11'd1541:   rom = 8'b00000000;    // 5
            11'd1542:   rom = 8'b00000000;    // 6
            11'd1543:   rom = 8'b00000000;    // 7
            11'd1544:   rom = 8'b00000000;    // 8
            11'd1545:   rom = 8'b00000000;    // 9
            11'd1546:   rom = 8'b00000000;    // a
            11'd1547:   rom = 8'b00000000;    // b
            11'd1548:   rom = 8'b00000000;    // c
            11'd1549:   rom = 8'b00000000;    // d
            11'd1550:   rom = 8'b00000000;    // e
            11'd1551:   rom = 8'b00000000;    // f
   // code x61
            11'd1552:   rom = 8'b00000000;    // 0
            11'd1553:   rom = 8'b00000000;    // 1
            11'd1554:   rom = 8'b00000000;    // 2
            11'd1555:   rom = 8'b00000000;    // 3
            11'd1556:   rom = 8'b00000000;    // 4
            11'd1557:   rom = 8'b01111000;    // 5  ****
            11'd1558:   rom = 8'b00001100;    // 6     **
            11'd1559:   rom = 8'b01111100;    // 7  *****
            11'd1560:   rom = 8'b11001100;    // 8 **  **
            11'd1561:   rom = 8'b11001100;    // 9 **  **
            11'd1562:   rom = 8'b11001100;    // a **  **
            11'd1563:   rom = 8'b01110110;    // b  *** **
            11'd1564:   rom = 8'b00000000;    // c
            11'd1565:   rom = 8'b00000000;    // d
            11'd1566:   rom = 8'b00000000;    // e
            11'd1567:   rom = 8'b00000000;    // f
   // code x62
            11'd1568:   rom = 8'b00000000;    // 0
            11'd1569:   rom = 8'b00000000;    // 1
            11'd1570:   rom = 8'b11100000;    // 2  ***
            11'd1571:   rom = 8'b01100000;    // 3   **
            11'd1572:   rom = 8'b01100000;    // 4   **
            11'd1573:   rom = 8'b01111000;    // 5   ****
            11'd1574:   rom = 8'b01101100;    // 6   ** **
            11'd1575:   rom = 8'b01100110;    // 7   **  **
            11'd1576:   rom = 8'b01100110;    // 8   **  **
            11'd1577:   rom = 8'b01100110;    // 9   **  **
            11'd1578:   rom = 8'b01100110;    // a   **  **
            11'd1579:   rom = 8'b01111100;    // b   *****
            11'd1580:   rom = 8'b00000000;    // c
            11'd1581:   rom = 8'b00000000;    // d
            11'd1582:   rom = 8'b00000000;    // e
            11'd1583:   rom = 8'b00000000;    // f
   // code x63
            11'd1584:   rom = 8'b00000000;    // 0
            11'd1585:   rom = 8'b00000000;    // 1
            11'd1586:   rom = 8'b00000000;    // 2
            11'd1587:   rom = 8'b00000000;    // 3
            11'd1588:   rom = 8'b00000000;    // 4
            11'd1589:   rom = 8'b01111100;    // 5  *****
            11'd1590:   rom = 8'b11000110;    // 6 **   **
            11'd1591:   rom = 8'b11000000;    // 7 **
            11'd1592:   rom = 8'b11000000;    // 8 **
            11'd1593:   rom = 8'b11000000;    // 9 **
            11'd1594:   rom = 8'b11000110;    // a **   **
            11'd1595:   rom = 8'b01111100;    // b  *****
            11'd1596:   rom = 8'b00000000;    // c
            11'd1597:   rom = 8'b00000000;    // d
            11'd1598:   rom = 8'b00000000;    // e
            11'd1599:   rom = 8'b00000000;    // f
   // code x64
            11'd1600:   rom = 8'b00000000;    // 0
            11'd1601:   rom = 8'b00000000;    // 1
            11'd1602:   rom = 8'b00011100;    // 2    ***
            11'd1603:   rom = 8'b00001100;    // 3     **
            11'd1604:   rom = 8'b00001100;    // 4     **
            11'd1605:   rom = 8'b00111100;    // 5   ****
            11'd1606:   rom = 8'b01101100;    // 6  ** **
            11'd1607:   rom = 8'b11001100;    // 7 **  **
            11'd1608:   rom = 8'b11001100;    // 8 **  **
            11'd1609:   rom = 8'b11001100;    // 9 **  **
            11'd1610:   rom = 8'b11001100;    // a **  **
            11'd1611:   rom = 8'b01110110;    // b  *** **
            11'd1612:   rom = 8'b00000000;    // c
            11'd1613:   rom = 8'b00000000;    // d
            11'd1614:   rom = 8'b00000000;    // e
            11'd1615:   rom = 8'b00000000;    // f
   // code x65
            11'd1616:   rom = 8'b00000000;    // 0
            11'd1617:   rom = 8'b00000000;    // 1
            11'd1618:   rom = 8'b00000000;    // 2
            11'd1619:   rom = 8'b00000000;    // 3
            11'd1620:   rom = 8'b00000000;    // 4
            11'd1621:   rom = 8'b01111100;    // 5  *****
            11'd1622:   rom = 8'b11000110;    // 6 **   **
            11'd1623:   rom = 8'b11111110;    // 7 *******
            11'd1624:   rom = 8'b11000000;    // 8 **
            11'd1625:   rom = 8'b11000000;    // 9 **
            11'd1626:   rom = 8'b11000110;    // a **   **
            11'd1627:   rom = 8'b01111100;    // b  *****
            11'd1628:   rom = 8'b00000000;    // c
            11'd1629:   rom = 8'b00000000;    // d
            11'd1630:   rom = 8'b00000000;    // e
            11'd1631:   rom = 8'b00000000;    // f
   // code x66
            11'd1632:   rom = 8'b00000000;    // 0
            11'd1633:   rom = 8'b00000000;    // 1
            11'd1634:   rom = 8'b00111000;    // 2   ***
            11'd1635:   rom = 8'b01101100;    // 3  ** **
            11'd1636:   rom = 8'b01100100;    // 4  **  *
            11'd1637:   rom = 8'b01100000;    // 5  **
            11'd1638:   rom = 8'b11110000;    // 6 ****
            11'd1639:   rom = 8'b01100000;    // 7  **
            11'd1640:   rom = 8'b01100000;    // 8  **
            11'd1641:   rom = 8'b01100000;    // 9  **
            11'd1642:   rom = 8'b01100000;    // a  **
            11'd1643:   rom = 8'b11110000;    // b ****
            11'd1644:   rom = 8'b00000000;    // c
            11'd1645:   rom = 8'b00000000;    // d
            11'd1646:   rom = 8'b00000000;    // e
            11'd1647:   rom = 8'b00000000;    // f
   // code x67
            11'd1648:   rom = 8'b00000000;    // 0
            11'd1649:   rom = 8'b00000000;    // 1
            11'd1650:   rom = 8'b00000000;    // 2
            11'd1651:   rom = 8'b00000000;    // 3
            11'd1652:   rom = 8'b00000000;    // 4
            11'd1653:   rom = 8'b01110110;    // 5  *** **
            11'd1654:   rom = 8'b11001100;    // 6 **  **
            11'd1655:   rom = 8'b11001100;    // 7 **  **
            11'd1656:   rom = 8'b11001100;    // 8 **  **
            11'd1657:   rom = 8'b11001100;    // 9 **  **
            11'd1658:   rom = 8'b11001100;    // a **  **
            11'd1659:   rom = 8'b01111100;    // b  *****
            11'd1660:   rom = 8'b00001100;    // c     **
            11'd1661:   rom = 8'b11001100;    // d **  **
            11'd1662:   rom = 8'b01111000;    // e  ****
            11'd1663:   rom = 8'b00000000;    // f
   // code x68
            11'd1664:   rom = 8'b00000000;    // 0
            11'd1665:   rom = 8'b00000000;    // 1
            11'd1666:   rom = 8'b11100000;    // 2 ***
            11'd1667:   rom = 8'b01100000;    // 3  **
            11'd1668:   rom = 8'b01100000;    // 4  **
            11'd1669:   rom = 8'b01101100;    // 5  ** **
            11'd1670:   rom = 8'b01110110;    // 6  *** **
            11'd1671:   rom = 8'b01100110;    // 7  **  **
            11'd1672:   rom = 8'b01100110;    // 8  **  **
            11'd1673:   rom = 8'b01100110;    // 9  **  **
            11'd1674:   rom = 8'b01100110;    // a  **  **
            11'd1675:   rom = 8'b11100110;    // b ***  **
            11'd1676:   rom = 8'b00000000;    // c
            11'd1677:   rom = 8'b00000000;    // d
            11'd1678:   rom = 8'b00000000;    // e
            11'd1679:   rom = 8'b00000000;    // f
   // code x69
            11'd1680:   rom = 8'b00000000;    // 0
            11'd1681:   rom = 8'b00000000;    // 1
            11'd1682:   rom = 8'b00011000;    // 2    **
            11'd1683:   rom = 8'b00011000;    // 3    **
            11'd1684:   rom = 8'b00000000;    // 4
            11'd1685:   rom = 8'b00111000;    // 5   ***
            11'd1686:   rom = 8'b00011000;    // 6    **
            11'd1687:   rom = 8'b00011000;    // 7    **
            11'd1688:   rom = 8'b00011000;    // 8    **
            11'd1689:   rom = 8'b00011000;    // 9    **
            11'd1690:   rom = 8'b00011000;    // a    **
            11'd1691:   rom = 8'b00111100;    // b   ****
            11'd1692:   rom = 8'b00000000;    // c
            11'd1693:   rom = 8'b00000000;    // d
            11'd1694:   rom = 8'b00000000;    // e
            11'd1695:   rom = 8'b00000000;    // f
   // code x6a
            11'd1696:   rom = 8'b00000000;    // 0
            11'd1697:   rom = 8'b00000000;    // 1
            11'd1698:   rom = 8'b00000110;    // 2      **
            11'd1699:   rom = 8'b00000110;    // 3      **
            11'd1700:   rom = 8'b00000000;    // 4
            11'd1701:   rom = 8'b00001110;    // 5     ***
            11'd1702:   rom = 8'b00000110;    // 6      **
            11'd1703:   rom = 8'b00000110;    // 7      **
            11'd1704:   rom = 8'b00000110;    // 8      **
            11'd1705:   rom = 8'b00000110;    // 9      **
            11'd1706:   rom = 8'b00000110;    // a      **
            11'd1707:   rom = 8'b00000110;    // b      **
            11'd1708:   rom = 8'b01100110;    // c  **  **
            11'd1709:   rom = 8'b01100110;    // d  **  **
            11'd1710:   rom = 8'b00111100;    // e   ****
            11'd1711:   rom = 8'b00000000;    // f
   // code x6b
            11'd1712:   rom = 8'b00000000;    // 0
            11'd1713:   rom = 8'b00000000;    // 1
            11'd1714:   rom = 8'b11100000;    // 2 ***
            11'd1715:   rom = 8'b01100000;    // 3  **
            11'd1716:   rom = 8'b01100000;    // 4  **
            11'd1717:   rom = 8'b01100110;    // 5  **  **
            11'd1718:   rom = 8'b01101100;    // 6  ** **
            11'd1719:   rom = 8'b01111000;    // 7  ****
            11'd1720:   rom = 8'b01111000;    // 8  ****
            11'd1721:   rom = 8'b01101100;    // 9  ** **
            11'd1722:   rom = 8'b01100110;    // a  **  **
            11'd1723:   rom = 8'b11100110;    // b ***  **
            11'd1724:   rom = 8'b00000000;    // c
            11'd1725:   rom = 8'b00000000;    // d
            11'd1726:   rom = 8'b00000000;    // e
            11'd1727:   rom = 8'b00000000;    // f
   // code x6c
            11'd1728:   rom = 8'b00000000;    // 0
            11'd1729:   rom = 8'b00000000;    // 1
            11'd1730:   rom = 8'b00111000;    // 2   ***
            11'd1731:   rom = 8'b00011000;    // 3    **
            11'd1732:   rom = 8'b00011000;    // 4    **
            11'd1733:   rom = 8'b00011000;    // 5    **
            11'd1734:   rom = 8'b00011000;    // 6    **
            11'd1735:   rom = 8'b00011000;    // 7    **
            11'd1736:   rom = 8'b00011000;    // 8    **
            11'd1737:   rom = 8'b00011000;    // 9    **
            11'd1738:   rom = 8'b00011000;    // a    **
            11'd1739:   rom = 8'b00111100;    // b   ****
            11'd1740:   rom = 8'b00000000;    // c
            11'd1741:   rom = 8'b00000000;    // d
            11'd1742:   rom = 8'b00000000;    // e
            11'd1743:   rom = 8'b00000000;    // f
   // code x6d
            11'd1744:   rom = 8'b00000000;    // 0
            11'd1745:   rom = 8'b00000000;    // 1
            11'd1746:   rom = 8'b00000000;    // 2
            11'd1747:   rom = 8'b00000000;    // 3
            11'd1748:   rom = 8'b00000000;    // 4
            11'd1749:   rom = 8'b11100110;    // 5 ***  **
            11'd1750:   rom = 8'b11111111;    // 6 ********
            11'd1751:   rom = 8'b11011011;    // 7 ** ** **
            11'd1752:   rom = 8'b11011011;    // 8 ** ** **
            11'd1753:   rom = 8'b11011011;    // 9 ** ** **
            11'd1754:   rom = 8'b11011011;    // a ** ** **
            11'd1755:   rom = 8'b11011011;    // b ** ** **
            11'd1756:   rom = 8'b00000000;    // c
            11'd1757:   rom = 8'b00000000;    // d
            11'd1758:   rom = 8'b00000000;    // e
            11'd1759:   rom = 8'b00000000;    // f
   // code x6e
            11'd1760:   rom = 8'b00000000;    // 0
            11'd1761:   rom = 8'b00000000;    // 1
            11'd1762:   rom = 8'b00000000;    // 2
            11'd1763:   rom = 8'b00000000;    // 3
            11'd1764:   rom = 8'b00000000;    // 4
            11'd1765:   rom = 8'b11011100;    // 5 ** ***
            11'd1766:   rom = 8'b01100110;    // 6  **  **
            11'd1767:   rom = 8'b01100110;    // 7  **  **
            11'd1768:   rom = 8'b01100110;    // 8  **  **
            11'd1769:   rom = 8'b01100110;    // 9  **  **
            11'd1770:   rom = 8'b01100110;    // a  **  **
            11'd1771:   rom = 8'b01100110;    // b  **  **
            11'd1772:   rom = 8'b00000000;    // c
            11'd1773:   rom = 8'b00000000;    // d
            11'd1774:   rom = 8'b00000000;    // e
            11'd1775:   rom = 8'b00000000;    // f
   // code x6f
            11'd1776:   rom = 8'b00000000;    // 0
            11'd1777:   rom = 8'b00000000;    // 1
            11'd1778:   rom = 8'b00000000;    // 2
            11'd1779:   rom = 8'b00000000;    // 3
            11'd1780:   rom = 8'b00000000;    // 4
            11'd1781:   rom = 8'b01111100;    // 5  *****
            11'd1782:   rom = 8'b11000110;    // 6 **   **
            11'd1783:   rom = 8'b11000110;    // 7 **   **
            11'd1784:   rom = 8'b11000110;    // 8 **   **
            11'd1785:   rom = 8'b11000110;    // 9 **   **
            11'd1786:   rom = 8'b11000110;    // a **   **
            11'd1787:   rom = 8'b01111100;    // b  *****
            11'd1788:   rom = 8'b00000000;    // c
            11'd1789:   rom = 8'b00000000;    // d
            11'd1790:   rom = 8'b00000000;    // e
            11'd1791:   rom = 8'b00000000;    // f
   // code x70
            11'd1792:   rom = 8'b00000000;    // 0
            11'd1793:   rom = 8'b00000000;    // 1
            11'd1794:   rom = 8'b00000000;    // 2
            11'd1795:   rom = 8'b00000000;    // 3
            11'd1796:   rom = 8'b00000000;    // 4
            11'd1797:   rom = 8'b11011100;    // 5 ** ***
            11'd1798:   rom = 8'b01100110;    // 6  **  **
            11'd1799:   rom = 8'b01100110;    // 7  **  **
            11'd1800:   rom = 8'b01100110;    // 8  **  **
            11'd1801:   rom = 8'b01100110;    // 9  **  **
            11'd1802:   rom = 8'b01100110;    // a  **  **
            11'd1803:   rom = 8'b01111100;    // b  *****
            11'd1804:   rom = 8'b01100000;    // c  **
            11'd1805:   rom = 8'b01100000;    // d  **
            11'd1806:   rom = 8'b11110000;    // e ****
            11'd1807:   rom = 8'b00000000;    // f
   // code x71
            11'd1808:   rom = 8'b00000000;    // 0
            11'd1809:   rom = 8'b00000000;    // 1
            11'd1810:   rom = 8'b00000000;    // 2
            11'd1811:   rom = 8'b00000000;    // 3
            11'd1812:   rom = 8'b00000000;    // 4
            11'd1813:   rom = 8'b01110110;    // 5  *** **
            11'd1814:   rom = 8'b11001100;    // 6 **  **
            11'd1815:   rom = 8'b11001100;    // 7 **  **
            11'd1816:   rom = 8'b11001100;    // 8 **  **
            11'd1817:   rom = 8'b11001100;    // 9 **  **
            11'd1818:   rom = 8'b11001100;    // a **  **
            11'd1819:   rom = 8'b01111100;    // b  *****
            11'd1820:   rom = 8'b00001100;    // c     **
            11'd1821:   rom = 8'b00001100;    // d     **
            11'd1822:   rom = 8'b00011110;    // e    ****
            11'd1823:   rom = 8'b00000000;    // f
   // code x72
            11'd1824:   rom = 8'b00000000;    // 0
            11'd1825:   rom = 8'b00000000;    // 1
            11'd1826:   rom = 8'b00000000;    // 2
            11'd1827:   rom = 8'b00000000;    // 3
            11'd1828:   rom = 8'b00000000;    // 4
            11'd1829:   rom = 8'b11011100;    // 5 ** ***
            11'd1830:   rom = 8'b01110110;    // 6  *** **
            11'd1831:   rom = 8'b01100110;    // 7  **  **
            11'd1832:   rom = 8'b01100000;    // 8  **
            11'd1833:   rom = 8'b01100000;    // 9  **
            11'd1834:   rom = 8'b01100000;    // a  **
            11'd1835:   rom = 8'b11110000;    // b ****
            11'd1836:   rom = 8'b00000000;    // c
            11'd1837:   rom = 8'b00000000;    // d
            11'd1838:   rom = 8'b00000000;    // e
            11'd1839:   rom = 8'b00000000;    // f
   // code x73
            11'd1840:   rom = 8'b00000000;    // 0
            11'd1841:   rom = 8'b00000000;    // 1
            11'd1842:   rom = 8'b00000000;    // 2
            11'd1843:   rom = 8'b00000000;    // 3
            11'd1844:   rom = 8'b00000000;    // 4
            11'd1845:   rom = 8'b01111100;    // 5  *****
            11'd1846:   rom = 8'b11000110;    // 6 **   **
            11'd1847:   rom = 8'b01100000;    // 7  **
            11'd1848:   rom = 8'b00111000;    // 8   ***
            11'd1849:   rom = 8'b00001100;    // 9     **
            11'd1850:   rom = 8'b11000110;    // a **   **
            11'd1851:   rom = 8'b01111100;    // b  *****
            11'd1852:   rom = 8'b00000000;    // c
            11'd1853:   rom = 8'b00000000;    // d
            11'd1854:   rom = 8'b00000000;    // e
            11'd1855:   rom = 8'b00000000;    // f
   // code x74
            11'd1856:   rom = 8'b00000000;    // 0
            11'd1857:   rom = 8'b00000000;    // 1
            11'd1858:   rom = 8'b00010000;    // 2    *
            11'd1859:   rom = 8'b00110000;    // 3   **
            11'd1860:   rom = 8'b00110000;    // 4   **
            11'd1861:   rom = 8'b11111100;    // 5 ******
            11'd1862:   rom = 8'b00110000;    // 6   **
            11'd1863:   rom = 8'b00110000;    // 7   **
            11'd1864:   rom = 8'b00110000;    // 8   **
            11'd1865:   rom = 8'b00110000;    // 9   **
            11'd1866:   rom = 8'b00110110;    // a   ** **
            11'd1867:   rom = 8'b00011100;    // b    ***
            11'd1868:   rom = 8'b00000000;    // c
            11'd1869:   rom = 8'b00000000;    // d
            11'd1870:   rom = 8'b00000000;    // e
            11'd1871:   rom = 8'b00000000;    // f
   // code x75
            11'd1872:   rom = 8'b00000000;    // 0
            11'd1873:   rom = 8'b00000000;    // 1
            11'd1874:   rom = 8'b00000000;    // 2
            11'd1875:   rom = 8'b00000000;    // 3
            11'd1876:   rom = 8'b00000000;    // 4
            11'd1877:   rom = 8'b11001100;    // 5 **  **
            11'd1878:   rom = 8'b11001100;    // 6 **  **
            11'd1879:   rom = 8'b11001100;    // 7 **  **
            11'd1880:   rom = 8'b11001100;    // 8 **  **
            11'd1881:   rom = 8'b11001100;    // 9 **  **
            11'd1882:   rom = 8'b11001100;    // a **  **
            11'd1883:   rom = 8'b01110110;    // b  *** **
            11'd1884:   rom = 8'b00000000;    // c
            11'd1885:   rom = 8'b00000000;    // d
            11'd1886:   rom = 8'b00000000;    // e
            11'd1887:   rom = 8'b00000000;    // f
   // code x76
            11'd1888:   rom = 8'b00000000;    // 0
            11'd1889:   rom = 8'b00000000;    // 1
            11'd1890:   rom = 8'b00000000;    // 2
            11'd1891:   rom = 8'b00000000;    // 3
            11'd1892:   rom = 8'b00000000;    // 4
            11'd1893:   rom = 8'b11000011;    // 5 **    **
            11'd1894:   rom = 8'b11000011;    // 6 **    **
            11'd1895:   rom = 8'b11000011;    // 7 **    **
            11'd1896:   rom = 8'b11000011;    // 8 **    **
            11'd1897:   rom = 8'b01100110;    // 9  **  **
            11'd1898:   rom = 8'b00111100;    // a   ****
            11'd1899:   rom = 8'b00011000;    // b    **
            11'd1900:   rom = 8'b00000000;    // c
            11'd1901:   rom = 8'b00000000;    // d
            11'd1902:   rom = 8'b00000000;    // e
            11'd1903:   rom = 8'b00000000;    // f
   // code x77
            11'd1904:   rom = 8'b00000000;    // 0
            11'd1905:   rom = 8'b00000000;    // 1
            11'd1906:   rom = 8'b00000000;    // 2
            11'd1907:   rom = 8'b00000000;    // 3
            11'd1908:   rom = 8'b00000000;    // 4
            11'd1909:   rom = 8'b11000011;    // 5 **    **
            11'd1910:   rom = 8'b11000011;    // 6 **    **
            11'd1911:   rom = 8'b11000011;    // 7 **    **
            11'd1912:   rom = 8'b11011011;    // 8 ** ** **
            11'd1913:   rom = 8'b11011011;    // 9 ** ** **
            11'd1914:   rom = 8'b11111111;    // a ********
            11'd1915:   rom = 8'b01100110;    // b  **  **
            11'd1916:   rom = 8'b00000000;    // c
            11'd1917:   rom = 8'b00000000;    // d
            11'd1918:   rom = 8'b00000000;    // e
            11'd1919:   rom = 8'b00000000;    // f
   // code x78
            11'd1920:   rom = 8'b00000000;    // 0
            11'd1921:   rom = 8'b00000000;    // 1
            11'd1922:   rom = 8'b00000000;    // 2
            11'd1923:   rom = 8'b00000000;    // 3
            11'd1924:   rom = 8'b00000000;    // 4
            11'd1925:   rom = 8'b11000011;    // 5 **    **
            11'd1926:   rom = 8'b01100110;    // 6  **  **
            11'd1927:   rom = 8'b00111100;    // 7   ****
            11'd1928:   rom = 8'b00011000;    // 8    **
            11'd1929:   rom = 8'b00111100;    // 9   ****
            11'd1930:   rom = 8'b01100110;    // a  **  **
            11'd1931:   rom = 8'b11000011;    // b **    **
            11'd1932:   rom = 8'b00000000;    // c
            11'd1933:   rom = 8'b00000000;    // d
            11'd1934:   rom = 8'b00000000;    // e
            11'd1935:   rom = 8'b00000000;    // f
   // code x79
            11'd1936:   rom = 8'b00000000;    // 0
            11'd1937:   rom = 8'b00000000;    // 1
            11'd1938:   rom = 8'b00000000;    // 2
            11'd1939:   rom = 8'b00000000;    // 3
            11'd1940:   rom = 8'b00000000;    // 4
            11'd1941:   rom = 8'b11000110;    // 5 **   **
            11'd1942:   rom = 8'b11000110;    // 6 **   **
            11'd1943:   rom = 8'b11000110;    // 7 **   **
            11'd1944:   rom = 8'b11000110;    // 8 **   **
            11'd1945:   rom = 8'b11000110;    // 9 **   **
            11'd1946:   rom = 8'b11000110;    // a **   **
            11'd1947:   rom = 8'b01111110;    // b  ******
            11'd1948:   rom = 8'b00000110;    // c      **
            11'd1949:   rom = 8'b00001100;    // d     **
            11'd1950:   rom = 8'b11111000;    // e *****
            11'd1951:   rom = 8'b00000000;    // f
   // code x7a
            11'd1952:   rom = 8'b00000000;    // 0
            11'd1953:   rom = 8'b00000000;    // 1
            11'd1954:   rom = 8'b00000000;    // 2
            11'd1955:   rom = 8'b00000000;    // 3
            11'd1956:   rom = 8'b00000000;    // 4
            11'd1957:   rom = 8'b11111110;    // 5 *******
            11'd1958:   rom = 8'b11001100;    // 6 **  **
            11'd1959:   rom = 8'b00011000;    // 7    **
            11'd1960:   rom = 8'b00110000;    // 8   **
            11'd1961:   rom = 8'b01100000;    // 9  **
            11'd1962:   rom = 8'b11000110;    // a **   **
            11'd1963:   rom = 8'b11111110;    // b *******
            11'd1964:   rom = 8'b00000000;    // c
            11'd1965:   rom = 8'b00000000;    // d
            11'd1966:   rom = 8'b00000000;    // e
            11'd1967:   rom = 8'b00000000;    // f
   // code x7b
            11'd1968:   rom = 8'b00000000;    // 0
            11'd1969:   rom = 8'b00000000;    // 1
            11'd1970:   rom = 8'b00001110;    // 2     ***
            11'd1971:   rom = 8'b00011000;    // 3    **
            11'd1972:   rom = 8'b00011000;    // 4    **
            11'd1973:   rom = 8'b00011000;    // 5    **
            11'd1974:   rom = 8'b01110000;    // 6  ***
            11'd1975:   rom = 8'b00011000;    // 7    **
            11'd1976:   rom = 8'b00011000;    // 8    **
            11'd1977:   rom = 8'b00011000;    // 9    **
            11'd1978:   rom = 8'b00011000;    // a    **
            11'd1979:   rom = 8'b00001110;    // b     ***
            11'd1980:   rom = 8'b00000000;    // c
            11'd1981:   rom = 8'b00000000;    // d
            11'd1982:   rom = 8'b00000000;    // e
            11'd1983:   rom = 8'b00000000;    // f
   // code x7c
            11'd1984:   rom = 8'b00000000;    // 0
            11'd1985:   rom = 8'b00000000;    // 1
            11'd1986:   rom = 8'b00011000;    // 2    **
            11'd1987:   rom = 8'b00011000;    // 3    **
            11'd1988:   rom = 8'b00011000;    // 4    **
            11'd1989:   rom = 8'b00011000;    // 5    **
            11'd1990:   rom = 8'b00000000;    // 6
            11'd1991:   rom = 8'b00011000;    // 7    **
            11'd1992:   rom = 8'b00011000;    // 8    **
            11'd1993:   rom = 8'b00011000;    // 9    **
            11'd1994:   rom = 8'b00011000;    // a    **
            11'd1995:   rom = 8'b00011000;    // b    **
            11'd1996:   rom = 8'b00000000;    // c
            11'd1997:   rom = 8'b00000000;    // d
            11'd1998:   rom = 8'b00000000;    // e
            11'd1999:   rom = 8'b00000000;    // f
   // code x7d
            11'd2000:   rom = 8'b00000000;    // 0
            11'd2001:   rom = 8'b00000000;    // 1
            11'd2002:   rom = 8'b01110000;    // 2  ***
            11'd2003:   rom = 8'b00011000;    // 3    **
            11'd2004:   rom = 8'b00011000;    // 4    **
            11'd2005:   rom = 8'b00011000;    // 5    **
            11'd2006:   rom = 8'b00001110;    // 6     ***
            11'd2007:   rom = 8'b00011000;    // 7    **
            11'd2008:   rom = 8'b00011000;    // 8    **
            11'd2009:   rom = 8'b00011000;    // 9    **
            11'd2010:   rom = 8'b00011000;    // a    **
            11'd2011:   rom = 8'b01110000;    // b  ***
            11'd2012:   rom = 8'b00000000;    // c
            11'd2013:   rom = 8'b00000000;    // d
            11'd2014:   rom = 8'b00000000;    // e
            11'd2015:   rom = 8'b00000000;    // f
   // code x7e
            11'd2016:   rom = 8'b00000000;    // 0
            11'd2017:   rom = 8'b00000000;    // 1
            11'd2018:   rom = 8'b01110110;    // 2  *** **
            11'd2019:   rom = 8'b11011100;    // 3 ** ***
            11'd2020:   rom = 8'b00000000;    // 4
            11'd2021:   rom = 8'b00000000;    // 5
            11'd2022:   rom = 8'b00000000;    // 6
            11'd2023:   rom = 8'b00000000;    // 7
            11'd2024:   rom = 8'b00000000;    // 8
            11'd2025:   rom = 8'b00000000;    // 9
            11'd2026:   rom = 8'b00000000;    // a
            11'd2027:   rom = 8'b00000000;    // b
            11'd2028:   rom = 8'b00000000;    // c
            11'd2029:   rom = 8'b00000000;    // d
            11'd2030:   rom = 8'b00000000;    // e
            11'd2031:   rom = 8'b00000000;    // f
   // code x7f
            11'd2032:   rom = 8'b00000000;    // 0
            11'd2033:   rom = 8'b00000000;    // 1
            11'd2034:   rom = 8'b00000000;    // 2
            11'd2035:   rom = 8'b00000000;    // 3
            11'd2036:   rom = 8'b00010000;    // 4    *
            11'd2037:   rom = 8'b00111000;    // 5   ***
            11'd2038:   rom = 8'b01101100;    // 6  ** **
            11'd2039:   rom = 8'b11000110;    // 7 **   **
            11'd2040:   rom = 8'b11000110;    // 8 **   **
            11'd2041:   rom = 8'b11000110;    // 9 **   **
            11'd2042:   rom = 8'b11111110;    // a *******
            11'd2043:   rom = 8'b00000000;    // b
            11'd2044:   rom = 8'b00000000;    // c
            11'd2045:   rom = 8'b00000000;    // d
            11'd2046:   rom = 8'b00000000;    // e
     endcase
	end
endmodule
